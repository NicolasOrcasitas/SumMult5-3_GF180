VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO suma_mult_TOP
  CLASS BLOCK ;
  FOREIGN suma_mult_TOP ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN X[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 310.800 0.000 311.360 4.000 ;
    END
  END X[0]
  PIN X[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 495.600 0.000 496.160 4.000 ;
    END
  END X[10]
  PIN X[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 0.000 514.640 4.000 ;
    END
  END X[11]
  PIN X[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.560 0.000 533.120 4.000 ;
    END
  END X[12]
  PIN X[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 0.000 551.600 4.000 ;
    END
  END X[13]
  PIN X[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 569.520 0.000 570.080 4.000 ;
    END
  END X[14]
  PIN X[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 0.000 588.560 4.000 ;
    END
  END X[15]
  PIN X[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 606.480 0.000 607.040 4.000 ;
    END
  END X[16]
  PIN X[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 0.000 625.520 4.000 ;
    END
  END X[17]
  PIN X[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 643.440 0.000 644.000 4.000 ;
    END
  END X[18]
  PIN X[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 0.000 662.480 4.000 ;
    END
  END X[19]
  PIN X[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 0.000 329.840 4.000 ;
    END
  END X[1]
  PIN X[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 680.400 0.000 680.960 4.000 ;
    END
  END X[20]
  PIN X[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 0.000 699.440 4.000 ;
    END
  END X[21]
  PIN X[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 717.360 0.000 717.920 4.000 ;
    END
  END X[22]
  PIN X[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 0.000 736.400 4.000 ;
    END
  END X[23]
  PIN X[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 754.320 0.000 754.880 4.000 ;
    END
  END X[24]
  PIN X[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 0.000 773.360 4.000 ;
    END
  END X[25]
  PIN X[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 791.280 0.000 791.840 4.000 ;
    END
  END X[26]
  PIN X[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 0.000 810.320 4.000 ;
    END
  END X[27]
  PIN X[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 828.240 0.000 828.800 4.000 ;
    END
  END X[28]
  PIN X[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 846.720 0.000 847.280 4.000 ;
    END
  END X[29]
  PIN X[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 347.760 0.000 348.320 4.000 ;
    END
  END X[2]
  PIN X[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 865.200 0.000 865.760 4.000 ;
    END
  END X[30]
  PIN X[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 0.000 884.240 4.000 ;
    END
  END X[31]
  PIN X[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END X[3]
  PIN X[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.720 0.000 385.280 4.000 ;
    END
  END X[4]
  PIN X[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 0.000 403.760 4.000 ;
    END
  END X[5]
  PIN X[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 421.680 0.000 422.240 4.000 ;
    END
  END X[6]
  PIN X[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 0.000 440.720 4.000 ;
    END
  END X[7]
  PIN X[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.640 0.000 459.200 4.000 ;
    END
  END X[8]
  PIN X[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 0.000 477.680 4.000 ;
    END
  END X[9]
  PIN b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 299.600 900.000 300.160 ;
    END
  END b
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 449.680 596.000 450.240 600.000 ;
    END
  END clk
  PIN n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.120 0.000 15.680 4.000 ;
    END
  END n[0]
  PIN n[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.920 0.000 200.480 4.000 ;
    END
  END n[10]
  PIN n[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END n[11]
  PIN n[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.880 0.000 237.440 4.000 ;
    END
  END n[12]
  PIN n[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END n[13]
  PIN n[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.840 0.000 274.400 4.000 ;
    END
  END n[14]
  PIN n[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 0.000 292.880 4.000 ;
    END
  END n[15]
  PIN n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END n[1]
  PIN n[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.080 0.000 52.640 4.000 ;
    END
  END n[2]
  PIN n[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END n[3]
  PIN n[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.040 0.000 89.600 4.000 ;
    END
  END n[4]
  PIN n[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END n[5]
  PIN n[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.000 0.000 126.560 4.000 ;
    END
  END n[6]
  PIN n[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END n[7]
  PIN n[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.960 0.000 163.520 4.000 ;
    END
  END n[8]
  PIN n[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 0.000 182.000 4.000 ;
    END
  END n[9]
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 299.600 4.000 300.160 ;
    END
  END start
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 584.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 893.200 584.380 ;
      LAYER Metal2 ;
        RECT 9.100 595.700 449.380 596.000 ;
        RECT 450.540 595.700 886.900 596.000 ;
        RECT 9.100 4.300 886.900 595.700 ;
        RECT 9.100 4.000 14.820 4.300 ;
        RECT 15.980 4.000 33.300 4.300 ;
        RECT 34.460 4.000 51.780 4.300 ;
        RECT 52.940 4.000 70.260 4.300 ;
        RECT 71.420 4.000 88.740 4.300 ;
        RECT 89.900 4.000 107.220 4.300 ;
        RECT 108.380 4.000 125.700 4.300 ;
        RECT 126.860 4.000 144.180 4.300 ;
        RECT 145.340 4.000 162.660 4.300 ;
        RECT 163.820 4.000 181.140 4.300 ;
        RECT 182.300 4.000 199.620 4.300 ;
        RECT 200.780 4.000 218.100 4.300 ;
        RECT 219.260 4.000 236.580 4.300 ;
        RECT 237.740 4.000 255.060 4.300 ;
        RECT 256.220 4.000 273.540 4.300 ;
        RECT 274.700 4.000 292.020 4.300 ;
        RECT 293.180 4.000 310.500 4.300 ;
        RECT 311.660 4.000 328.980 4.300 ;
        RECT 330.140 4.000 347.460 4.300 ;
        RECT 348.620 4.000 365.940 4.300 ;
        RECT 367.100 4.000 384.420 4.300 ;
        RECT 385.580 4.000 402.900 4.300 ;
        RECT 404.060 4.000 421.380 4.300 ;
        RECT 422.540 4.000 439.860 4.300 ;
        RECT 441.020 4.000 458.340 4.300 ;
        RECT 459.500 4.000 476.820 4.300 ;
        RECT 477.980 4.000 495.300 4.300 ;
        RECT 496.460 4.000 513.780 4.300 ;
        RECT 514.940 4.000 532.260 4.300 ;
        RECT 533.420 4.000 550.740 4.300 ;
        RECT 551.900 4.000 569.220 4.300 ;
        RECT 570.380 4.000 587.700 4.300 ;
        RECT 588.860 4.000 606.180 4.300 ;
        RECT 607.340 4.000 624.660 4.300 ;
        RECT 625.820 4.000 643.140 4.300 ;
        RECT 644.300 4.000 661.620 4.300 ;
        RECT 662.780 4.000 680.100 4.300 ;
        RECT 681.260 4.000 698.580 4.300 ;
        RECT 699.740 4.000 717.060 4.300 ;
        RECT 718.220 4.000 735.540 4.300 ;
        RECT 736.700 4.000 754.020 4.300 ;
        RECT 755.180 4.000 772.500 4.300 ;
        RECT 773.660 4.000 790.980 4.300 ;
        RECT 792.140 4.000 809.460 4.300 ;
        RECT 810.620 4.000 827.940 4.300 ;
        RECT 829.100 4.000 846.420 4.300 ;
        RECT 847.580 4.000 864.900 4.300 ;
        RECT 866.060 4.000 883.380 4.300 ;
        RECT 884.540 4.000 886.900 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 300.460 896.000 584.220 ;
        RECT 4.300 299.300 895.700 300.460 ;
        RECT 4.000 11.900 896.000 299.300 ;
      LAYER Metal4 ;
        RECT 159.180 28.090 175.540 198.150 ;
        RECT 177.740 28.090 252.340 198.150 ;
        RECT 254.540 28.090 329.140 198.150 ;
        RECT 331.340 28.090 405.940 198.150 ;
        RECT 408.140 28.090 482.740 198.150 ;
        RECT 484.940 28.090 559.540 198.150 ;
        RECT 561.740 28.090 636.340 198.150 ;
        RECT 638.540 28.090 686.980 198.150 ;
  END
END suma_mult_TOP
END LIBRARY

