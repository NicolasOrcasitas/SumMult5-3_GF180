// This is the unpowered netlist.
module suma_mult_TOP (b,
    clk,
    start,
    X,
    n);
 output b;
 input clk;
 input start;
 output [31:0] X;
 input [15:0] n;

 wire \Control_Unit.C[0] ;
 wire \Control_Unit.C[10] ;
 wire \Control_Unit.C[11] ;
 wire \Control_Unit.C[12] ;
 wire \Control_Unit.C[13] ;
 wire \Control_Unit.C[14] ;
 wire \Control_Unit.C[15] ;
 wire \Control_Unit.C[16] ;
 wire \Control_Unit.C[17] ;
 wire \Control_Unit.C[18] ;
 wire \Control_Unit.C[19] ;
 wire \Control_Unit.C[1] ;
 wire \Control_Unit.C[20] ;
 wire \Control_Unit.C[21] ;
 wire \Control_Unit.C[22] ;
 wire \Control_Unit.C[23] ;
 wire \Control_Unit.C[24] ;
 wire \Control_Unit.C[25] ;
 wire \Control_Unit.C[26] ;
 wire \Control_Unit.C[27] ;
 wire \Control_Unit.C[28] ;
 wire \Control_Unit.C[29] ;
 wire \Control_Unit.C[2] ;
 wire \Control_Unit.C[30] ;
 wire \Control_Unit.C[31] ;
 wire \Control_Unit.C[3] ;
 wire \Control_Unit.C[4] ;
 wire \Control_Unit.C[5] ;
 wire \Control_Unit.C[6] ;
 wire \Control_Unit.C[7] ;
 wire \Control_Unit.C[8] ;
 wire \Control_Unit.C[9] ;
 wire \Control_Unit.Mc ;
 wire \Control_Unit.Mq ;
 wire \Control_Unit.Mt ;
 wire \Control_Unit.Mx ;
 wire \Control_Unit.Q[0] ;
 wire \Control_Unit.Q[10] ;
 wire \Control_Unit.Q[11] ;
 wire \Control_Unit.Q[12] ;
 wire \Control_Unit.Q[13] ;
 wire \Control_Unit.Q[14] ;
 wire \Control_Unit.Q[15] ;
 wire \Control_Unit.Q[16] ;
 wire \Control_Unit.Q[17] ;
 wire \Control_Unit.Q[18] ;
 wire \Control_Unit.Q[19] ;
 wire \Control_Unit.Q[1] ;
 wire \Control_Unit.Q[20] ;
 wire \Control_Unit.Q[21] ;
 wire \Control_Unit.Q[22] ;
 wire \Control_Unit.Q[23] ;
 wire \Control_Unit.Q[24] ;
 wire \Control_Unit.Q[25] ;
 wire \Control_Unit.Q[26] ;
 wire \Control_Unit.Q[27] ;
 wire \Control_Unit.Q[28] ;
 wire \Control_Unit.Q[29] ;
 wire \Control_Unit.Q[2] ;
 wire \Control_Unit.Q[30] ;
 wire \Control_Unit.Q[31] ;
 wire \Control_Unit.Q[3] ;
 wire \Control_Unit.Q[4] ;
 wire \Control_Unit.Q[5] ;
 wire \Control_Unit.Q[6] ;
 wire \Control_Unit.Q[7] ;
 wire \Control_Unit.Q[8] ;
 wire \Control_Unit.Q[9] ;
 wire \Control_Unit.Rc ;
 wire \Control_Unit.Rcont ;
 wire \Control_Unit.Rx ;
 wire \Control_Unit.T[0] ;
 wire \Control_Unit.T[10] ;
 wire \Control_Unit.T[11] ;
 wire \Control_Unit.T[12] ;
 wire \Control_Unit.T[13] ;
 wire \Control_Unit.T[14] ;
 wire \Control_Unit.T[15] ;
 wire \Control_Unit.T[16] ;
 wire \Control_Unit.T[17] ;
 wire \Control_Unit.T[18] ;
 wire \Control_Unit.T[19] ;
 wire \Control_Unit.T[1] ;
 wire \Control_Unit.T[20] ;
 wire \Control_Unit.T[21] ;
 wire \Control_Unit.T[22] ;
 wire \Control_Unit.T[23] ;
 wire \Control_Unit.T[24] ;
 wire \Control_Unit.T[25] ;
 wire \Control_Unit.T[26] ;
 wire \Control_Unit.T[27] ;
 wire \Control_Unit.T[28] ;
 wire \Control_Unit.T[29] ;
 wire \Control_Unit.T[2] ;
 wire \Control_Unit.T[30] ;
 wire \Control_Unit.T[31] ;
 wire \Control_Unit.T[3] ;
 wire \Control_Unit.T[4] ;
 wire \Control_Unit.T[5] ;
 wire \Control_Unit.T[6] ;
 wire \Control_Unit.T[7] ;
 wire \Control_Unit.T[8] ;
 wire \Control_Unit.T[9] ;
 wire \Control_Unit.cont[0] ;
 wire \Control_Unit.cont[10] ;
 wire \Control_Unit.cont[11] ;
 wire \Control_Unit.cont[12] ;
 wire \Control_Unit.cont[13] ;
 wire \Control_Unit.cont[14] ;
 wire \Control_Unit.cont[15] ;
 wire \Control_Unit.cont[1] ;
 wire \Control_Unit.cont[2] ;
 wire \Control_Unit.cont[3] ;
 wire \Control_Unit.cont[4] ;
 wire \Control_Unit.cont[5] ;
 wire \Control_Unit.cont[6] ;
 wire \Control_Unit.cont[7] ;
 wire \Control_Unit.cont[8] ;
 wire \Control_Unit.cont[9] ;
 wire \Control_Unit.futuro[0] ;
 wire \Control_Unit.futuro[1] ;
 wire \Control_Unit.futuro[2] ;
 wire \Control_Unit.presente[0] ;
 wire \Control_Unit.presente[1] ;
 wire \Control_Unit.presente[2] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;

 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2335_ (.I(\Control_Unit.presente[2] ),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2336_ (.I(\Control_Unit.presente[1] ),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2337_ (.A1(_1673_),
    .A2(_1674_),
    .A3(\Control_Unit.presente[0] ),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2338_ (.I(_1675_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2339_ (.I(\Control_Unit.presente[0] ),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2340_ (.I(\Control_Unit.presente[1] ),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2341_ (.A1(_1673_),
    .A2(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2342_ (.I(_1678_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2343_ (.A1(_1676_),
    .A2(_1679_),
    .B(_1675_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2344_ (.I(\Control_Unit.presente[2] ),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2345_ (.I(\Control_Unit.presente[0] ),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2346_ (.A1(_1680_),
    .A2(_1681_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2347_ (.A1(\Control_Unit.presente[2] ),
    .A2(_1674_),
    .A3(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2348_ (.A1(_1675_),
    .A2(_1682_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2349_ (.I(\Control_Unit.presente[0] ),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2350_ (.A1(\Control_Unit.presente[2] ),
    .A2(_1677_),
    .A3(_1683_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2351_ (.A1(_1677_),
    .A2(_1683_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2352_ (.A1(_1673_),
    .A2(_1685_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2353_ (.I(_1686_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2354_ (.A1(_1684_),
    .A2(_0007_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2355_ (.A1(_1675_),
    .A2(_1679_),
    .A3(_1682_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2356_ (.A1(_1680_),
    .A2(_1676_),
    .B(_1684_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2357_ (.A1(_1679_),
    .A2(_1682_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2358_ (.I(net10),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2359_ (.I(net9),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2360_ (.I(net15),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2361_ (.I(_1689_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2362_ (.I(net14),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2363_ (.I(net13),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2364_ (.I(net12),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2365_ (.A1(_1690_),
    .A2(_1691_),
    .A3(_1692_),
    .A4(_1693_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2366_ (.I(net4),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2367_ (.I(net3),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2368_ (.I(net17),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2369_ (.I(net16),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2370_ (.A1(_1695_),
    .A2(_1696_),
    .A3(_1697_),
    .A4(_1698_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2371_ (.I(net5),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2372_ (.A1(net8),
    .A2(net7),
    .A3(net6),
    .A4(_1700_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2373_ (.A1(_1694_),
    .A2(_1699_),
    .A3(_1701_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2374_ (.I(net11),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2375_ (.A1(_1687_),
    .A2(_1688_),
    .B(_1702_),
    .C(_1703_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2376_ (.I(_1704_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2377_ (.I(\Control_Unit.cont[15] ),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2378_ (.I(_1706_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2379_ (.I(_1707_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2380_ (.I(\Control_Unit.cont[14] ),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2381_ (.I(_1709_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2382_ (.I(\Control_Unit.cont[12] ),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2383_ (.I(\Control_Unit.cont[13] ),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2384_ (.I(\Control_Unit.cont[11] ),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2385_ (.I(\Control_Unit.cont[8] ),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2386_ (.I(\Control_Unit.cont[9] ),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2387_ (.I(\Control_Unit.cont[10] ),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2388_ (.I(\Control_Unit.cont[6] ),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2389_ (.I(\Control_Unit.cont[7] ),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2390_ (.A1(\Control_Unit.cont[3] ),
    .A2(\Control_Unit.cont[2] ),
    .A3(\Control_Unit.cont[1] ),
    .A4(\Control_Unit.cont[0] ),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2391_ (.A1(\Control_Unit.cont[4] ),
    .A2(\Control_Unit.cont[5] ),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2392_ (.A1(_1717_),
    .A2(_1718_),
    .A3(_1719_),
    .A4(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2393_ (.I(_1721_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2394_ (.A1(_1714_),
    .A2(_1715_),
    .A3(_1716_),
    .A4(_1722_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2395_ (.A1(_1713_),
    .A2(_1723_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2396_ (.A1(_1711_),
    .A2(_1712_),
    .A3(_1724_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2397_ (.A1(_1710_),
    .A2(_1725_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2398_ (.I(_1726_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2399_ (.I(\Control_Unit.cont[15] ),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2400_ (.A1(_1710_),
    .A2(_1725_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2401_ (.A1(_1728_),
    .A2(_1729_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2402_ (.A1(_1727_),
    .A2(_1730_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2403_ (.A1(_1708_),
    .A2(_1727_),
    .B(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2404_ (.I(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2405_ (.I(\Control_Unit.cont[14] ),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2406_ (.I(\Control_Unit.cont[13] ),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2407_ (.I(\Control_Unit.cont[12] ),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2408_ (.A1(_1736_),
    .A2(_1724_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2409_ (.A1(_1735_),
    .A2(_1737_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2410_ (.A1(_1734_),
    .A2(_1738_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2411_ (.A1(_1726_),
    .A2(_1738_),
    .B(_1739_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2412_ (.I(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2413_ (.A1(_1713_),
    .A2(_1723_),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2414_ (.A1(\Control_Unit.cont[12] ),
    .A2(_1724_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2415_ (.A1(_1736_),
    .A2(_1742_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2416_ (.A1(_1742_),
    .A2(_1743_),
    .B(_1744_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2417_ (.I(\Control_Unit.cont[9] ),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2418_ (.A1(\Control_Unit.cont[8] ),
    .A2(_1722_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2419_ (.A1(_1746_),
    .A2(_1747_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2420_ (.I(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2421_ (.I(_1749_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2422_ (.I(_1750_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2423_ (.I(_1714_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2424_ (.A1(_1752_),
    .A2(_1722_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2425_ (.I(_1753_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2426_ (.I(_1754_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2427_ (.A1(_1751_),
    .A2(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2428_ (.I(\Control_Unit.cont[8] ),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2429_ (.A1(_1757_),
    .A2(_1722_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2430_ (.I(_1714_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2431_ (.I(\Control_Unit.cont[7] ),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2432_ (.A1(_1717_),
    .A2(_1719_),
    .A3(_1720_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2433_ (.A1(_1760_),
    .A2(_1761_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2434_ (.I0(_1758_),
    .I1(_1759_),
    .S(_1762_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2435_ (.I(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2436_ (.I(_1760_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2437_ (.I(_1765_),
    .Z(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2438_ (.I(_1766_),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2439_ (.I(_1767_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2440_ (.I(\Control_Unit.cont[3] ),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2441_ (.I(\Control_Unit.cont[0] ),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2442_ (.A1(_1769_),
    .A2(\Control_Unit.cont[2] ),
    .A3(\Control_Unit.cont[1] ),
    .A4(_1770_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2443_ (.I(_1771_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2444_ (.I(\Control_Unit.cont[4] ),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2445_ (.I(\Control_Unit.cont[5] ),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2446_ (.A1(_1773_),
    .A2(_1774_),
    .Z(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2447_ (.I(\Control_Unit.cont[6] ),
    .Z(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2448_ (.A1(_1772_),
    .A2(_1775_),
    .B(_1776_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2449_ (.A1(_1761_),
    .A2(_1777_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2450_ (.I(_1778_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2451_ (.I(_1779_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2452_ (.I(_1762_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2453_ (.A1(_1781_),
    .A2(_1778_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2454_ (.I(_1774_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2455_ (.I(_1783_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2456_ (.I(_1773_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2457_ (.A1(_1785_),
    .A2(_1772_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2458_ (.I(_1786_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2459_ (.A1(_1784_),
    .A2(_1787_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2460_ (.A1(_1772_),
    .A2(_1775_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2461_ (.A1(_1785_),
    .A2(_1719_),
    .B(_1784_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2462_ (.A1(_1773_),
    .A2(_1771_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2463_ (.I(_1791_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2464_ (.I(_1792_),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2465_ (.A1(_1789_),
    .A2(_1790_),
    .B(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2466_ (.I(\Control_Unit.cont[2] ),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2467_ (.I(_1795_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2468_ (.I(_1796_),
    .Z(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2469_ (.I(_1797_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2470_ (.I(_1798_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2471_ (.I(\Control_Unit.cont[1] ),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2472_ (.I(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2473_ (.I(_1801_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2474_ (.I(_1770_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2475_ (.I(_1803_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2476_ (.A1(_1802_),
    .A2(_1804_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2477_ (.I(_1805_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2478_ (.I(_1802_),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2479_ (.I(_1807_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2480_ (.I(_1808_),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2481_ (.I(_1770_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2482_ (.I(_1810_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2483_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2484_ (.I(_1812_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2485_ (.I(_1813_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2486_ (.A1(_1795_),
    .A2(_1800_),
    .A3(_1810_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2487_ (.I(_1815_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2488_ (.A1(_1801_),
    .A2(_1811_),
    .B(_1796_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2489_ (.A1(_1809_),
    .A2(_1814_),
    .B1(_1816_),
    .B2(_1817_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2490_ (.I(_1769_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2491_ (.I(_1819_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2492_ (.I(_1820_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2493_ (.I(_1821_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2494_ (.A1(_1799_),
    .A2(_1806_),
    .B1(_1818_),
    .B2(_1822_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2495_ (.I(\Control_Unit.cont[4] ),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2496_ (.I(_1824_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2497_ (.I(_1825_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2498_ (.A1(_1819_),
    .A2(_1815_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2499_ (.I(_1827_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2500_ (.I0(_1787_),
    .I1(_1826_),
    .S(_1828_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2501_ (.A1(_1788_),
    .A2(_1794_),
    .A3(_1823_),
    .A4(_1829_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2502_ (.I(_1774_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2503_ (.I(_1831_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2504_ (.A1(_1832_),
    .A2(_1791_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2505_ (.I(_1827_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2506_ (.I(_1834_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(_1826_),
    .A2(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2508_ (.A1(_1833_),
    .A2(_1836_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2509_ (.I(_1776_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2510_ (.I(_1838_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2511_ (.A1(_1839_),
    .A2(_1789_),
    .A3(_1790_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2512_ (.A1(_1824_),
    .A2(_1772_),
    .B(_1774_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2513_ (.I(_1841_),
    .Z(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2514_ (.A1(_1719_),
    .A2(_1720_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2515_ (.I(_1843_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2516_ (.A1(_1761_),
    .A2(_1777_),
    .B1(_1842_),
    .B2(_1844_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2517_ (.A1(_1840_),
    .A2(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2518_ (.A1(_1830_),
    .A2(_1837_),
    .B(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2519_ (.I(_1717_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2520_ (.A1(_1848_),
    .A2(_1844_),
    .A3(_1842_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2521_ (.A1(_1768_),
    .A2(_1780_),
    .B1(_1782_),
    .B2(_1847_),
    .C(_1849_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2522_ (.A1(_1756_),
    .A2(_1764_),
    .A3(_1850_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2523_ (.I(_1715_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2524_ (.A1(_1852_),
    .A2(_1753_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2525_ (.A1(_1759_),
    .A2(_1781_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2526_ (.A1(_1853_),
    .A2(_1854_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2527_ (.I(_1742_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2528_ (.I(_1716_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2529_ (.A1(\Control_Unit.cont[8] ),
    .A2(\Control_Unit.cont[9] ),
    .A3(_1721_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2530_ (.A1(_1857_),
    .A2(_1858_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2531_ (.I(_1859_),
    .Z(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2532_ (.A1(_1856_),
    .A2(_1860_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2533_ (.A1(_1716_),
    .A2(_1748_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2534_ (.A1(\Control_Unit.cont[10] ),
    .A2(_1858_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2535_ (.A1(\Control_Unit.cont[9] ),
    .A2(_1747_),
    .Z(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2536_ (.A1(_1863_),
    .A2(_1864_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2537_ (.A1(_1862_),
    .A2(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2538_ (.A1(_1851_),
    .A2(_1855_),
    .B(_1861_),
    .C(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2539_ (.I(\Control_Unit.cont[11] ),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2540_ (.A1(_1868_),
    .A2(_1859_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2541_ (.A1(_1869_),
    .A2(_1862_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2542_ (.A1(_1867_),
    .A2(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2543_ (.A1(_1745_),
    .A2(_1871_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2544_ (.I(_1738_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2545_ (.I(_1873_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2546_ (.I(_1743_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2547_ (.I(_1875_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2548_ (.I(_1876_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2549_ (.A1(_1874_),
    .A2(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2550_ (.I(_1712_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2551_ (.I(_1879_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2552_ (.I(_1880_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2553_ (.I(_1881_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2554_ (.A1(_1882_),
    .A2(_1877_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2555_ (.A1(_1872_),
    .A2(_1878_),
    .B(_1744_),
    .C(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2556_ (.A1(_1741_),
    .A2(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2557_ (.A1(_1739_),
    .A2(_1885_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2558_ (.A1(_1733_),
    .A2(_1886_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2559_ (.I(net6),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2560_ (.I(_1735_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2561_ (.I0(_1873_),
    .I1(_1889_),
    .S(_1875_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2562_ (.A1(_1744_),
    .A2(_1872_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2563_ (.A1(_1890_),
    .A2(_1891_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2564_ (.A1(_1851_),
    .A2(_1855_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2565_ (.A1(_1866_),
    .A2(_1893_),
    .B(_1862_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2566_ (.A1(_1856_),
    .A2(_1860_),
    .B(_1869_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2567_ (.A1(_1894_),
    .A2(_1895_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2568_ (.A1(_1866_),
    .A2(_1893_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2569_ (.A1(_1764_),
    .A2(_1850_),
    .B(_1854_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2570_ (.A1(_1748_),
    .A2(_1753_),
    .B(_1853_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2571_ (.A1(_1898_),
    .A2(_1899_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2572_ (.A1(_1697_),
    .A2(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2573_ (.A1(_1764_),
    .A2(_1850_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2574_ (.A1(_1849_),
    .A2(_1847_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2575_ (.I0(_1762_),
    .I1(_1718_),
    .S(_1778_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2576_ (.A1(_1903_),
    .A2(_1904_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2577_ (.A1(_1689_),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2578_ (.A1(_1830_),
    .A2(_1837_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2579_ (.A1(_1846_),
    .A2(_1907_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2580_ (.I(net12),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2581_ (.I(_1785_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2582_ (.I0(_1792_),
    .I1(_1910_),
    .S(_1827_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2583_ (.A1(_1823_),
    .A2(_1911_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2584_ (.I(_1828_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2585_ (.I(_1769_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2586_ (.I(_1914_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2587_ (.I(_1915_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2588_ (.A1(_1816_),
    .A2(_1817_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2589_ (.I(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2590_ (.I0(_1913_),
    .I1(_1916_),
    .S(_1918_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2591_ (.I(_1799_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2592_ (.I(_1814_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2593_ (.A1(_1809_),
    .A2(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2594_ (.A1(_1920_),
    .A2(_1806_),
    .B(_1922_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2595_ (.A1(_1919_),
    .A2(_1923_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2596_ (.I(_1807_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2597_ (.I(_1925_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2598_ (.I(_1926_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2599_ (.I(_1921_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2600_ (.A1(_1927_),
    .A2(net9),
    .B1(net2),
    .B2(_1928_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2601_ (.A1(_1921_),
    .A2(net2),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2602_ (.A1(_1927_),
    .A2(net9),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2603_ (.A1(_1929_),
    .A2(_1930_),
    .B(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2604_ (.I(_1797_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2605_ (.I(_1933_),
    .Z(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2606_ (.A1(_1934_),
    .A2(_1928_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2607_ (.A1(net10),
    .A2(_1932_),
    .B(_1935_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2608_ (.I(net10),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2609_ (.A1(_1937_),
    .A2(_1932_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2610_ (.A1(net11),
    .A2(_1924_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2611_ (.A1(_1936_),
    .A2(_1938_),
    .B(_1939_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2612_ (.A1(_1909_),
    .A2(_1912_),
    .B1(_1924_),
    .B2(net11),
    .C(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2613_ (.A1(_1823_),
    .A2(_1829_),
    .B(_1836_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2614_ (.A1(_1843_),
    .A2(_1841_),
    .B(_1786_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2615_ (.A1(_1833_),
    .A2(_1943_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2616_ (.A1(_1942_),
    .A2(_1944_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2617_ (.A1(net13),
    .A2(_1945_),
    .B1(_1912_),
    .B2(_1909_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2618_ (.A1(_1691_),
    .A2(_1908_),
    .B1(_1945_),
    .B2(net13),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2619_ (.A1(_1941_),
    .A2(_1946_),
    .B(_1947_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2620_ (.A1(_1689_),
    .A2(_1905_),
    .B1(_1908_),
    .B2(_1691_),
    .C(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2621_ (.A1(net16),
    .A2(_1902_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2622_ (.A1(_1906_),
    .A2(_1949_),
    .B(_1950_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2623_ (.A1(net17),
    .A2(_1900_),
    .B1(_1902_),
    .B2(_1698_),
    .C(_1951_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2624_ (.A1(net3),
    .A2(_1897_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2625_ (.A1(_1901_),
    .A2(_1952_),
    .B(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2626_ (.A1(net4),
    .A2(_1896_),
    .B1(_1897_),
    .B2(_1696_),
    .C(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2627_ (.A1(_1745_),
    .A2(_1871_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2628_ (.A1(_1872_),
    .A2(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2629_ (.A1(net5),
    .A2(_1957_),
    .B1(_1896_),
    .B2(net4),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2630_ (.A1(net5),
    .A2(_1957_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2631_ (.A1(_1888_),
    .A2(_1892_),
    .B1(_1955_),
    .B2(_1958_),
    .C(_1959_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2632_ (.A1(_1740_),
    .A2(_1884_),
    .Z(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2633_ (.A1(net7),
    .A2(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2634_ (.A1(_1888_),
    .A2(_1892_),
    .B(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2635_ (.I(net7),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2636_ (.A1(net8),
    .A2(_1887_),
    .B1(_1960_),
    .B2(_1963_),
    .C1(_1961_),
    .C2(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2637_ (.I(_1708_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2638_ (.I(_1966_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2639_ (.A1(_1967_),
    .A2(_1729_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2640_ (.A1(_1968_),
    .A2(_1739_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2641_ (.I(net8),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2642_ (.A1(_1731_),
    .A2(_1885_),
    .B1(_1887_),
    .B2(_1970_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2643_ (.A1(_1965_),
    .A2(_1969_),
    .A3(_1971_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2644_ (.A1(_1676_),
    .A2(_1678_),
    .A3(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2645_ (.A1(_1705_),
    .A2(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2646_ (.A1(net18),
    .A2(_1684_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2647_ (.I(\Control_Unit.C[25] ),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2648_ (.I(\Control_Unit.C[24] ),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2649_ (.I(\Control_Unit.C[27] ),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2650_ (.I(\Control_Unit.C[26] ),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2651_ (.A1(_1976_),
    .A2(_1977_),
    .A3(_1978_),
    .A4(_1979_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2652_ (.I(\Control_Unit.C[21] ),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2653_ (.I(_1981_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2654_ (.I(\Control_Unit.C[20] ),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2655_ (.I(\Control_Unit.C[23] ),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2656_ (.I(\Control_Unit.C[22] ),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2657_ (.A1(_1982_),
    .A2(_1983_),
    .A3(_1984_),
    .A4(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2658_ (.I(\Control_Unit.C[17] ),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2659_ (.I(_1987_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2660_ (.I(\Control_Unit.C[16] ),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2661_ (.I(\Control_Unit.C[19] ),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2662_ (.I(_1990_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2663_ (.I(\Control_Unit.C[18] ),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2664_ (.I(_1992_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2665_ (.A1(_1988_),
    .A2(_1989_),
    .A3(_1991_),
    .A4(_1993_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2666_ (.I(\Control_Unit.C[29] ),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2667_ (.I(\Control_Unit.C[28] ),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2668_ (.I(\Control_Unit.C[30] ),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2669_ (.A1(_1995_),
    .A2(_1996_),
    .A3(\Control_Unit.C[31] ),
    .A4(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2670_ (.A1(_1986_),
    .A2(_1994_),
    .A3(_1998_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2671_ (.I(\Control_Unit.C[9] ),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2672_ (.I(\Control_Unit.C[8] ),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2673_ (.I(\Control_Unit.C[11] ),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2674_ (.I(_2002_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2675_ (.I(\Control_Unit.C[10] ),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2676_ (.A1(_2000_),
    .A2(_2001_),
    .A3(_2003_),
    .A4(_2004_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2677_ (.I(\Control_Unit.C[5] ),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2678_ (.I(_2006_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2679_ (.I(\Control_Unit.C[4] ),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2680_ (.I(_2008_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2681_ (.I(\Control_Unit.C[7] ),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2682_ (.I(\Control_Unit.C[6] ),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2683_ (.A1(_2007_),
    .A2(_2009_),
    .A3(_2010_),
    .A4(_2011_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2684_ (.I(\Control_Unit.C[1] ),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2685_ (.I(\Control_Unit.C[0] ),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2686_ (.I(\Control_Unit.C[3] ),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2687_ (.I(\Control_Unit.C[2] ),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2688_ (.A1(_2013_),
    .A2(_2014_),
    .A3(_2015_),
    .A4(_2016_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2689_ (.I(\Control_Unit.C[13] ),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2690_ (.I(\Control_Unit.C[12] ),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2691_ (.I(\Control_Unit.C[15] ),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2692_ (.I(\Control_Unit.C[14] ),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2693_ (.A1(_2018_),
    .A2(_2019_),
    .A3(_2020_),
    .A4(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2694_ (.A1(_2012_),
    .A2(_2017_),
    .A3(_2022_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2695_ (.A1(_1980_),
    .A2(_1999_),
    .A3(_2005_),
    .A4(_2023_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2696_ (.A1(_1680_),
    .A2(_1674_),
    .A3(_1683_),
    .A4(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2697_ (.I(_1734_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2698_ (.I(_2026_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2699_ (.A1(_2027_),
    .A2(_1876_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2700_ (.I(_2028_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2701_ (.I(_1856_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2702_ (.A1(_1880_),
    .A2(_2030_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2703_ (.A1(_1727_),
    .A2(_1876_),
    .B(_2028_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2704_ (.A1(_2031_),
    .A2(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2705_ (.A1(_1873_),
    .A2(_2030_),
    .B(_2031_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2706_ (.I(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2707_ (.I(_1868_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2708_ (.I(_2036_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2709_ (.A1(_2037_),
    .A2(_1749_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2710_ (.I(_2038_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2711_ (.I(_1860_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2712_ (.I(_1711_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2713_ (.A1(_2041_),
    .A2(_2040_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2714_ (.A1(_1875_),
    .A2(_2040_),
    .B(_2042_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2715_ (.A1(_2039_),
    .A2(_2043_),
    .B(_2042_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2716_ (.I(_1856_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2717_ (.I(\Control_Unit.cont[10] ),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2718_ (.I(_2046_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2719_ (.A1(_2047_),
    .A2(_1754_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2720_ (.A1(_2040_),
    .A2(_1755_),
    .B(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2721_ (.I(_1852_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2722_ (.I(_1781_),
    .Z(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2723_ (.A1(_2050_),
    .A2(_2051_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2724_ (.A1(_2049_),
    .A2(_2052_),
    .B(_2048_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2725_ (.A1(_2045_),
    .A2(_1751_),
    .B(_2039_),
    .C(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2726_ (.I(_2050_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2727_ (.I(_2051_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2728_ (.A1(_1750_),
    .A2(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2729_ (.A1(_2055_),
    .A2(_2056_),
    .B(_2057_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2730_ (.I(_1757_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2731_ (.I(_2059_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2732_ (.I(_1778_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2733_ (.A1(_1755_),
    .A2(_1780_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2734_ (.A1(_1844_),
    .A2(_1842_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2735_ (.I(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2736_ (.A1(_1767_),
    .A2(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2737_ (.I(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2738_ (.I(_1717_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2739_ (.I(_1787_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2740_ (.A1(_2067_),
    .A2(_2068_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2741_ (.I(_1832_),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2742_ (.A1(_2070_),
    .A2(_1835_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2743_ (.A1(_1910_),
    .A2(_1816_),
    .A3(_1817_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2744_ (.I(_1820_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2745_ (.A1(_2073_),
    .A2(_1805_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2746_ (.A1(_1934_),
    .A2(_1812_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2747_ (.A1(_1828_),
    .A2(_1806_),
    .B(_2075_),
    .C(_2074_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2748_ (.A1(_1793_),
    .A2(_1918_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2749_ (.A1(_2074_),
    .A2(_2076_),
    .B(_2072_),
    .C(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2750_ (.A1(_2064_),
    .A2(_1835_),
    .B1(_2072_),
    .B2(_2078_),
    .C(_2071_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2751_ (.A1(_1779_),
    .A2(_1787_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2752_ (.A1(_2071_),
    .A2(_2079_),
    .B(_2080_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2753_ (.I(_2064_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2754_ (.A1(_2066_),
    .A2(_2069_),
    .A3(_2081_),
    .B1(_2082_),
    .B2(_2056_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2755_ (.A1(_2060_),
    .A2(_2061_),
    .B1(_2062_),
    .B2(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2756_ (.A1(_2049_),
    .A2(_2052_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2757_ (.A1(_2030_),
    .A2(_1750_),
    .B(_2038_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2758_ (.A1(_2086_),
    .A2(_2048_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2759_ (.A1(_2058_),
    .A2(_2084_),
    .A3(_2085_),
    .A4(_2087_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2760_ (.A1(_2039_),
    .A2(_2043_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2761_ (.A1(_2054_),
    .A2(_2088_),
    .B(_2089_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2762_ (.A1(_2034_),
    .A2(_2042_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2763_ (.A1(_2035_),
    .A2(_2044_),
    .B1(_2090_),
    .B2(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2764_ (.A1(_2033_),
    .A2(_2092_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2765_ (.A1(_2031_),
    .A2(_2032_),
    .B(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2766_ (.A1(_1966_),
    .A2(_1874_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2767_ (.A1(_1730_),
    .A2(_1874_),
    .B(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2768_ (.A1(_2029_),
    .A2(_2094_),
    .A3(_2096_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2769_ (.A1(_2033_),
    .A2(_2092_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2770_ (.A1(_2093_),
    .A2(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2771_ (.A1(_2039_),
    .A2(_2043_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2772_ (.A1(_2100_),
    .A2(_2090_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2773_ (.A1(_2091_),
    .A2(_2101_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2774_ (.A1(net7),
    .A2(_2099_),
    .B1(_2102_),
    .B2(net6),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2775_ (.I(_2103_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2776_ (.A1(_2058_),
    .A2(_2084_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2777_ (.A1(_2052_),
    .A2(_2105_),
    .B(_2049_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2778_ (.A1(_2106_),
    .A2(_2087_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2779_ (.A1(_2105_),
    .A2(_2085_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2780_ (.A1(net3),
    .A2(_2108_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2781_ (.A1(_2058_),
    .A2(_2084_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2782_ (.I(_1759_),
    .Z(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2783_ (.I(_2111_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2784_ (.A1(_2112_),
    .A2(_1780_),
    .B(_2062_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2785_ (.A1(_2113_),
    .A2(_2083_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2786_ (.A1(net17),
    .A2(_2110_),
    .B1(_2114_),
    .B2(net16),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2787_ (.I(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2788_ (.A1(_2069_),
    .A2(_2081_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2789_ (.I(_2051_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2790_ (.A1(_2118_),
    .A2(_2082_),
    .B(_2065_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2791_ (.A1(_2117_),
    .A2(_2119_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2792_ (.A1(net16),
    .A2(_2114_),
    .B1(_2120_),
    .B2(_1689_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2793_ (.A1(net15),
    .A2(_2120_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2794_ (.I(net14),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2795_ (.A1(_2080_),
    .A2(_2071_),
    .A3(_2079_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2796_ (.A1(_2081_),
    .A2(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2797_ (.A1(_2123_),
    .A2(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2798_ (.A1(_2082_),
    .A2(_1913_),
    .B(_2071_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2799_ (.A1(_2072_),
    .A2(_2078_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2800_ (.A1(_2127_),
    .A2(_2128_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2801_ (.I(_2129_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2802_ (.A1(_1691_),
    .A2(_2081_),
    .A3(_2124_),
    .B1(_2130_),
    .B2(net13),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2803_ (.A1(_2126_),
    .A2(_2131_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2804_ (.I(_1918_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2805_ (.A1(_2074_),
    .A2(_2076_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2806_ (.A1(_2068_),
    .A2(_2133_),
    .A3(_2134_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2807_ (.A1(_1692_),
    .A2(_2130_),
    .B1(_2135_),
    .B2(_1909_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2808_ (.A1(_1909_),
    .A2(_2135_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2809_ (.A1(_1913_),
    .A2(_1806_),
    .B(_2074_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2810_ (.A1(_2075_),
    .A2(_2138_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2811_ (.A1(_1703_),
    .A2(_2139_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2812_ (.I(net11),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2813_ (.A1(_1928_),
    .A2(_2133_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2814_ (.A1(_2141_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(_1937_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2815_ (.A1(_1808_),
    .A2(_1813_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2816_ (.I(_2144_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2817_ (.A1(_1688_),
    .A2(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2818_ (.A1(_1688_),
    .A2(_2145_),
    .B1(_2142_),
    .B2(_1937_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2819_ (.I(_2147_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2820_ (.A1(_1930_),
    .A2(_2143_),
    .A3(_2146_),
    .A4(_2148_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2821_ (.A1(_2137_),
    .A2(_2140_),
    .A3(_2149_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2822_ (.A1(_2132_),
    .A2(_2136_),
    .A3(_2150_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2823_ (.A1(_2121_),
    .A2(_2122_),
    .A3(_2151_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2824_ (.I(_1928_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2825_ (.A1(_2153_),
    .A2(net2),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2826_ (.A1(_2154_),
    .A2(_2146_),
    .B(_2147_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2827_ (.A1(_1703_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(_1687_),
    .C(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2828_ (.A1(_2137_),
    .A2(_2140_),
    .A3(_2156_),
    .B(_2136_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2829_ (.A1(_2132_),
    .A2(_2157_),
    .B(_2122_),
    .C(_2126_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2830_ (.A1(_2121_),
    .A2(_2158_),
    .B(_2115_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2831_ (.A1(_1697_),
    .A2(_2110_),
    .B1(_2116_),
    .B2(_2152_),
    .C(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2832_ (.A1(net3),
    .A2(_2108_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2833_ (.A1(_2109_),
    .A2(_2160_),
    .B(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2834_ (.A1(_1695_),
    .A2(_2107_),
    .B(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2835_ (.A1(_2054_),
    .A2(_2088_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2836_ (.A1(_2164_),
    .A2(_2089_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2837_ (.A1(_1700_),
    .A2(_2165_),
    .B1(_2107_),
    .B2(_1695_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2838_ (.A1(net6),
    .A2(_2102_),
    .B1(_2165_),
    .B2(_1700_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2839_ (.A1(_2163_),
    .A2(_2166_),
    .B(_2167_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2840_ (.A1(net8),
    .A2(_2097_),
    .B1(_2104_),
    .B2(_2168_),
    .C1(_2099_),
    .C2(_1964_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2841_ (.A1(_2029_),
    .A2(_2096_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2842_ (.A1(_2029_),
    .A2(_2096_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2843_ (.A1(_2094_),
    .A2(_2170_),
    .B(_2171_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2844_ (.I(_1874_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2845_ (.I(_1727_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2846_ (.A1(_1967_),
    .A2(_2173_),
    .B(_2174_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2847_ (.I(_2027_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2848_ (.I(_2176_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2849_ (.A1(_2177_),
    .A2(_1966_),
    .B1(_1733_),
    .B2(_2173_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2850_ (.A1(_2174_),
    .A2(_2173_),
    .B(_2178_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2851_ (.A1(_2172_),
    .A2(_2179_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2852_ (.A1(_2172_),
    .A2(_2175_),
    .B(_2180_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2853_ (.A1(_1970_),
    .A2(_2097_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2854_ (.A1(_2177_),
    .A2(_1967_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2855_ (.A1(_1967_),
    .A2(_2174_),
    .B1(_2183_),
    .B2(_1725_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2856_ (.A1(_2169_),
    .A2(_2181_),
    .A3(_2182_),
    .A4(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2857_ (.A1(_1680_),
    .A2(_1685_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2858_ (.A1(_1702_),
    .A2(_2185_),
    .B(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2859_ (.A1(_1974_),
    .A2(_1975_),
    .A3(_2025_),
    .A4(_2187_),
    .ZN(\Control_Unit.futuro[0] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2860_ (.A1(_1881_),
    .A2(_1876_),
    .B1(_1890_),
    .B2(_2030_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2861_ (.A1(_1740_),
    .A2(_1875_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2862_ (.A1(_2188_),
    .A2(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2863_ (.I(_2045_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2864_ (.A1(_2188_),
    .A2(_2189_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2865_ (.A1(_2191_),
    .A2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2866_ (.A1(_2176_),
    .A2(_1877_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2867_ (.A1(_1890_),
    .A2(_2029_),
    .A3(_2194_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2868_ (.A1(_1732_),
    .A2(_1873_),
    .A3(_2195_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2869_ (.A1(_2190_),
    .A2(_2193_),
    .B(_2196_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2870_ (.A1(_2190_),
    .A2(_2193_),
    .A3(_2196_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2871_ (.A1(_2197_),
    .A2(_2198_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2872_ (.A1(_2045_),
    .A2(_2192_),
    .Z(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2873_ (.A1(_1745_),
    .A2(_1863_),
    .B(_1744_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2874_ (.A1(_2045_),
    .A2(_1890_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2875_ (.A1(_2201_),
    .A2(_2202_),
    .Z(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2876_ (.A1(_2201_),
    .A2(_2202_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2877_ (.A1(_2040_),
    .A2(_2203_),
    .B(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2878_ (.A1(_2200_),
    .A2(_2205_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2879_ (.A1(_2200_),
    .A2(_2205_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2880_ (.I(_2047_),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2881_ (.A1(_2208_),
    .A2(_1750_),
    .B1(_1865_),
    .B2(_1754_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2882_ (.A1(_1749_),
    .A2(_1895_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2883_ (.A1(_2209_),
    .A2(_2210_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2884_ (.A1(_2209_),
    .A2(_2210_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2885_ (.A1(_1758_),
    .A2(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2886_ (.A1(_1861_),
    .A2(_1864_),
    .B(_1869_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2887_ (.A1(_1745_),
    .A2(_1860_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2888_ (.A1(_2214_),
    .A2(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2889_ (.A1(_1751_),
    .A2(_2216_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2890_ (.A1(_2211_),
    .A2(_2213_),
    .B(_2217_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2891_ (.A1(_2217_),
    .A2(_2211_),
    .A3(_2213_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2892_ (.A1(_2218_),
    .A2(_2219_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2893_ (.A1(_1749_),
    .A2(_1754_),
    .B(_1853_),
    .C(_2051_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2894_ (.A1(_1853_),
    .A2(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2895_ (.A1(_1866_),
    .A2(_1753_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2896_ (.I(_2223_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2897_ (.A1(_2222_),
    .A2(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2898_ (.A1(_2222_),
    .A2(_2223_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2899_ (.A1(_2118_),
    .A2(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2900_ (.A1(_1755_),
    .A2(_2212_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2901_ (.A1(_2225_),
    .A2(_2227_),
    .B(_2228_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2902_ (.A1(_2118_),
    .A2(_2226_),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2903_ (.A1(_1764_),
    .A2(_2061_),
    .B(_1854_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2904_ (.I(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2905_ (.A1(_1781_),
    .A2(_1899_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2906_ (.A1(_2232_),
    .A2(_2233_),
    .Z(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2907_ (.A1(_2232_),
    .A2(_2233_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2908_ (.A1(_2061_),
    .A2(_2234_),
    .B(_2235_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2909_ (.A1(_2227_),
    .A2(_2230_),
    .A3(_2236_),
    .Z(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2910_ (.A1(_1845_),
    .A2(_1792_),
    .B(_1849_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2911_ (.A1(_2063_),
    .A2(_1904_),
    .A3(_2238_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2912_ (.A1(_1793_),
    .A2(_2239_),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2913_ (.A1(_1840_),
    .A2(_1845_),
    .A3(_1792_),
    .Z(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2914_ (.A1(_1840_),
    .A2(_1845_),
    .B(_1793_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2915_ (.A1(_1943_),
    .A2(_1834_),
    .B(_1788_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2916_ (.A1(_2241_),
    .A2(_2242_),
    .B(_2243_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2917_ (.A1(_2241_),
    .A2(_2243_),
    .A3(_2242_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2918_ (.A1(_1913_),
    .A2(_2244_),
    .B(_2245_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2919_ (.A1(_2240_),
    .A2(_2246_),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2920_ (.A1(_1916_),
    .A2(_1933_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2921_ (.A1(_1821_),
    .A2(_1917_),
    .B1(_1805_),
    .B2(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2922_ (.A1(_1918_),
    .A2(_1829_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2923_ (.A1(_2249_),
    .A2(_2250_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2924_ (.A1(_1917_),
    .A2(_1911_),
    .A3(_2249_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2925_ (.A1(_2145_),
    .A2(_2252_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2926_ (.A1(_2251_),
    .A2(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2927_ (.I(_1825_),
    .Z(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2928_ (.A1(_2255_),
    .A2(_1834_),
    .B1(_1917_),
    .B2(_1911_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2929_ (.A1(_1834_),
    .A2(_1944_),
    .A3(_2256_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2930_ (.A1(_2133_),
    .A2(_2257_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2931_ (.A1(_2254_),
    .A2(_2258_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2932_ (.A1(_1916_),
    .A2(_1934_),
    .A3(_1809_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2933_ (.A1(_1927_),
    .A2(_1919_),
    .B(_1921_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2934_ (.A1(_2144_),
    .A2(_2252_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2935_ (.A1(_2260_),
    .A2(_2261_),
    .A3(_2262_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2936_ (.A1(_2254_),
    .A2(_2258_),
    .B(_2263_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2937_ (.I(_1828_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2938_ (.A1(_2241_),
    .A2(_2242_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2939_ (.A1(_2265_),
    .A2(_2243_),
    .A3(_2266_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2940_ (.A1(_1788_),
    .A2(_1794_),
    .A3(_2265_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2941_ (.A1(_1833_),
    .A2(_1943_),
    .B(_1835_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2942_ (.A1(_2268_),
    .A2(_2256_),
    .A3(_2269_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2943_ (.A1(_2133_),
    .A2(_2257_),
    .B(_2270_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2944_ (.A1(_2267_),
    .A2(_2271_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2945_ (.A1(_2247_),
    .A2(_2259_),
    .A3(_2264_),
    .A4(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2946_ (.I(_1822_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2947_ (.A1(_2274_),
    .A2(_1920_),
    .A3(_1922_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2948_ (.A1(_1829_),
    .A2(_2275_),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2949_ (.A1(_2240_),
    .A2(_2246_),
    .B1(_2276_),
    .B2(_1944_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2950_ (.A1(_2240_),
    .A2(_2246_),
    .B(_2267_),
    .C(_2271_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2951_ (.A1(_2277_),
    .A2(_2278_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2952_ (.A1(_1766_),
    .A2(_1779_),
    .B1(_1782_),
    .B2(_2063_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2953_ (.A1(_1763_),
    .A2(_1779_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2954_ (.A1(_2063_),
    .A2(_2280_),
    .A3(_2281_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2955_ (.I(_2282_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2956_ (.A1(_2064_),
    .A2(_1904_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2957_ (.A1(_2238_),
    .A2(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2958_ (.A1(_2068_),
    .A2(_2239_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2959_ (.A1(_2285_),
    .A2(_2286_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2960_ (.A1(_2283_),
    .A2(_2287_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2961_ (.A1(_1780_),
    .A2(_2231_),
    .A3(_2233_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2962_ (.A1(_2280_),
    .A2(_2281_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2963_ (.A1(_2280_),
    .A2(_2281_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2964_ (.A1(_2082_),
    .A2(_2290_),
    .B(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2965_ (.A1(_2289_),
    .A2(_2292_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2966_ (.A1(_2273_),
    .A2(_2279_),
    .B(_2288_),
    .C(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2967_ (.A1(_2289_),
    .A2(_2292_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2968_ (.A1(_2283_),
    .A2(_2287_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2969_ (.A1(_2289_),
    .A2(_2292_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2970_ (.A1(_2295_),
    .A2(_2296_),
    .B(_2297_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2971_ (.A1(_2056_),
    .A2(_2226_),
    .A3(_2236_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2972_ (.A1(_2294_),
    .A2(_2298_),
    .B(_2299_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2973_ (.A1(_2225_),
    .A2(_2227_),
    .A3(_2228_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2974_ (.A1(_2229_),
    .A2(_2237_),
    .A3(_2300_),
    .B(_2301_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2975_ (.A1(_2220_),
    .A2(_2302_),
    .B(_2218_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2976_ (.A1(_1863_),
    .A2(_2201_),
    .A3(_2202_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2977_ (.I(_2215_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2978_ (.A1(_2214_),
    .A2(_2305_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2979_ (.A1(_1751_),
    .A2(_2216_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2980_ (.A1(_2304_),
    .A2(_2306_),
    .A3(_2307_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2981_ (.A1(_2306_),
    .A2(_2307_),
    .B(_2304_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2982_ (.A1(_2303_),
    .A2(_2308_),
    .B(_2309_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2983_ (.A1(_2207_),
    .A2(_2310_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2984_ (.A1(_2206_),
    .A2(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2985_ (.A1(_2199_),
    .A2(_2312_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2986_ (.A1(_2207_),
    .A2(_2310_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2987_ (.I(_2308_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2988_ (.A1(_2309_),
    .A2(_2315_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2989_ (.A1(_2303_),
    .A2(_2316_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2990_ (.A1(_2237_),
    .A2(_2300_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2991_ (.A1(_2225_),
    .A2(_2227_),
    .A3(_2228_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2992_ (.A1(_2229_),
    .A2(_2319_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2993_ (.A1(_2318_),
    .A2(_2320_),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2994_ (.A1(_2294_),
    .A2(_2298_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2995_ (.A1(_2299_),
    .A2(_2322_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2996_ (.A1(net4),
    .A2(_2321_),
    .B1(_2323_),
    .B2(_1696_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2997_ (.I(_1697_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2998_ (.A1(_2247_),
    .A2(_2259_),
    .A3(_2264_),
    .A4(_2272_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2999_ (.A1(_2277_),
    .A2(_2278_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3000_ (.A1(_2282_),
    .A2(_2287_),
    .Z(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3001_ (.A1(_2326_),
    .A2(_2327_),
    .B(_2328_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3002_ (.A1(_2296_),
    .A2(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3003_ (.A1(_2330_),
    .A2(_2293_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3004_ (.A1(_2273_),
    .A2(_2279_),
    .A3(_2288_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3005_ (.A1(_2329_),
    .A2(_2332_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3006_ (.A1(_1698_),
    .A2(_2333_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3007_ (.A1(_2325_),
    .A2(_2331_),
    .B(_2334_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3008_ (.A1(_2267_),
    .A2(_2271_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3009_ (.A1(_2267_),
    .A2(_2271_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3010_ (.A1(_0154_),
    .A2(_0155_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3011_ (.A1(_1944_),
    .A2(_2276_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3012_ (.A1(_2259_),
    .A2(_2264_),
    .B(_0157_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3013_ (.A1(_0156_),
    .A2(_0158_),
    .B(_0154_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3014_ (.A1(_2247_),
    .A2(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3015_ (.A1(_0156_),
    .A2(_0158_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3016_ (.A1(_2123_),
    .A2(_0161_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3017_ (.A1(_1690_),
    .A2(_0160_),
    .B(_0162_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3018_ (.A1(_2263_),
    .A2(_2275_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3019_ (.A1(_2254_),
    .A2(_2258_),
    .A3(_0164_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3020_ (.A1(_1692_),
    .A2(_0165_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3021_ (.A1(_2260_),
    .A2(_2261_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3022_ (.A1(_0167_),
    .A2(_2262_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3023_ (.A1(_2275_),
    .A2(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3024_ (.A1(_2276_),
    .A2(_0169_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3025_ (.A1(_1692_),
    .A2(_0165_),
    .B1(_0170_),
    .B2(_1693_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3026_ (.A1(_1931_),
    .A2(_1930_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3027_ (.A1(_2274_),
    .A2(_2141_),
    .B1(_1937_),
    .B2(_1920_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3028_ (.A1(_2274_),
    .A2(_2141_),
    .B1(_1687_),
    .B2(_1920_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3029_ (.A1(_1927_),
    .A2(_1688_),
    .B(_0174_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3030_ (.A1(_0172_),
    .A2(_0173_),
    .A3(_0175_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3031_ (.A1(_1693_),
    .A2(_0170_),
    .B(_0171_),
    .C(_0176_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3032_ (.A1(_2123_),
    .A2(_0161_),
    .B(_0166_),
    .C(_0177_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3033_ (.A1(_1698_),
    .A2(_2333_),
    .B1(_0160_),
    .B2(_1690_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3034_ (.A1(_2274_),
    .A2(_2141_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3035_ (.A1(_0180_),
    .A2(_0174_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3036_ (.A1(_1929_),
    .A2(_1931_),
    .B(_0173_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3037_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_0170_),
    .B2(_1693_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3038_ (.A1(_2123_),
    .A2(_0161_),
    .B1(_0171_),
    .B2(_0183_),
    .C(_0166_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3039_ (.A1(_1690_),
    .A2(_0160_),
    .B(_0162_),
    .C(_0184_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3040_ (.A1(_0163_),
    .A2(_0178_),
    .B(_0179_),
    .C(_0185_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3041_ (.A1(_2325_),
    .A2(_2331_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3042_ (.A1(_1696_),
    .A2(_2323_),
    .B1(_0153_),
    .B2(_0186_),
    .C(_0187_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3043_ (.A1(_2220_),
    .A2(_2302_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3044_ (.A1(net5),
    .A2(_0189_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3045_ (.A1(_1695_),
    .A2(_2321_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3046_ (.A1(_2324_),
    .A2(_0188_),
    .B(_0190_),
    .C(_0191_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3047_ (.A1(_1700_),
    .A2(_0189_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3048_ (.A1(_1888_),
    .A2(_2317_),
    .B(_0193_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3049_ (.A1(_1964_),
    .A2(_2314_),
    .B1(_0192_),
    .B2(_0194_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3050_ (.A1(_1888_),
    .A2(_2317_),
    .B(_0195_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3051_ (.A1(_1970_),
    .A2(_2313_),
    .B1(_2314_),
    .B2(_1964_),
    .C(_0196_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3052_ (.A1(_1970_),
    .A2(_2313_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3053_ (.A1(_2199_),
    .A2(_2311_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3054_ (.A1(_1889_),
    .A2(_1737_),
    .A3(_2183_),
    .A4(_2197_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3055_ (.A1(_2190_),
    .A2(_2193_),
    .A3(_2196_),
    .B(_2206_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3056_ (.A1(_0199_),
    .A2(_0200_),
    .A3(_0201_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3057_ (.I(_1682_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3058_ (.A1(_0197_),
    .A2(_0198_),
    .A3(_0202_),
    .B(_0203_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3059_ (.A1(_1703_),
    .A2(_1687_),
    .A3(_1702_),
    .B(_0152_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3060_ (.I(_1702_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3061_ (.A1(_0206_),
    .A2(_2185_),
    .B(_2186_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3062_ (.A1(_1683_),
    .A2(_1678_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3063_ (.A1(_1704_),
    .A2(_1972_),
    .B(_0208_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3064_ (.A1(_2025_),
    .A2(_0209_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3065_ (.A1(_0204_),
    .A2(_0205_),
    .A3(_0207_),
    .A4(_0210_),
    .ZN(\Control_Unit.futuro[1] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3066_ (.A1(_1676_),
    .A2(_2024_),
    .B(_1673_),
    .C(_1677_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3067_ (.A1(_1973_),
    .A2(_0211_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3068_ (.A1(_1681_),
    .A2(_1679_),
    .A3(_2185_),
    .B(_0212_),
    .ZN(\Control_Unit.futuro[2] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3069_ (.I(\Control_Unit.T[11] ),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3070_ (.A1(_2208_),
    .A2(_0213_),
    .A3(_2037_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3071_ (.I(_1857_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3072_ (.I(\Control_Unit.T[10] ),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3073_ (.A1(_2055_),
    .A2(_0216_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3074_ (.A1(_2055_),
    .A2(_0216_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3075_ (.A1(_0215_),
    .A2(_0217_),
    .B(_0218_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3076_ (.A1(_0214_),
    .A2(_0219_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3077_ (.I(_0220_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3078_ (.I(_2208_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3079_ (.A1(_2050_),
    .A2(_0216_),
    .A3(_0222_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3080_ (.I(_1746_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3081_ (.I(\Control_Unit.T[9] ),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3082_ (.A1(_2112_),
    .A2(_0225_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3083_ (.A1(_2112_),
    .A2(_0225_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3084_ (.A1(_0224_),
    .A2(_0226_),
    .B(_0227_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3085_ (.A1(_0223_),
    .A2(_0228_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3086_ (.A1(_2111_),
    .A2(\Control_Unit.T[9] ),
    .A3(_2050_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3087_ (.I(\Control_Unit.T[8] ),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3088_ (.A1(_1768_),
    .A2(_0231_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3089_ (.A1(_1768_),
    .A2(_0231_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3090_ (.A1(_2060_),
    .A2(_0232_),
    .B(_0233_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3091_ (.A1(_0230_),
    .A2(_0234_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3092_ (.I(_0235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3093_ (.A1(_1767_),
    .A2(\Control_Unit.T[8] ),
    .A3(_2111_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3094_ (.I(_1718_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3095_ (.I(_1839_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3096_ (.I(\Control_Unit.T[7] ),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3097_ (.A1(_0239_),
    .A2(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3098_ (.A1(_0239_),
    .A2(_0240_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3099_ (.A1(_0238_),
    .A2(_0241_),
    .B(_0242_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3100_ (.A1(_0237_),
    .A2(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3101_ (.I(_1832_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3102_ (.I(\Control_Unit.T[6] ),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3103_ (.A1(_0245_),
    .A2(_0246_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3104_ (.A1(_2070_),
    .A2(_0246_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3105_ (.A1(_0239_),
    .A2(_0248_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3106_ (.A1(_1848_),
    .A2(\Control_Unit.T[7] ),
    .A3(_1767_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3107_ (.A1(_0247_),
    .A2(_0249_),
    .B(_0250_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3108_ (.A1(_2067_),
    .A2(_0248_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3109_ (.A1(\Control_Unit.T[5] ),
    .A2(_2255_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3110_ (.I(\Control_Unit.T[5] ),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3111_ (.A1(_0254_),
    .A2(_1826_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3112_ (.A1(_0245_),
    .A2(_0253_),
    .B(_0255_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3113_ (.A1(_0252_),
    .A2(_0256_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3114_ (.A1(_0250_),
    .A2(_0247_),
    .A3(_0249_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3115_ (.A1(_0251_),
    .A2(_0257_),
    .B(_0258_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3116_ (.I(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3117_ (.A1(_0252_),
    .A2(_0256_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3118_ (.I(\Control_Unit.T[4] ),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3119_ (.I(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3120_ (.A1(_0262_),
    .A2(_2073_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3121_ (.A1(_1826_),
    .A2(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3122_ (.A1(_0263_),
    .A2(_1916_),
    .B(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3123_ (.A1(_0245_),
    .A2(_0253_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3124_ (.A1(_0266_),
    .A2(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3125_ (.I(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3126_ (.I(\Control_Unit.T[3] ),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3127_ (.A1(_1799_),
    .A2(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3128_ (.A1(_1798_),
    .A2(_0270_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3129_ (.A1(_1822_),
    .A2(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3130_ (.A1(_0271_),
    .A2(_0273_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3131_ (.A1(_2255_),
    .A2(_0264_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3132_ (.A1(_0274_),
    .A2(_0275_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3133_ (.I(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3134_ (.I(\Control_Unit.T[0] ),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3135_ (.A1(_1812_),
    .A2(\Control_Unit.T[1] ),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3136_ (.A1(_1925_),
    .A2(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3137_ (.A1(_1814_),
    .A2(_0278_),
    .A3(_0280_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3138_ (.I(_1801_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3139_ (.A1(_1933_),
    .A2(_0282_),
    .A3(\Control_Unit.T[2] ),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3140_ (.A1(_1812_),
    .A2(\Control_Unit.T[1] ),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3141_ (.A1(_1925_),
    .A2(_0279_),
    .B(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3142_ (.A1(_0283_),
    .A2(_0285_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3143_ (.A1(_0283_),
    .A2(_0285_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3144_ (.A1(_0281_),
    .A2(_0286_),
    .B(_0287_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3145_ (.A1(_1821_),
    .A2(_0272_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3146_ (.I(\Control_Unit.T[2] ),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3147_ (.A1(_1925_),
    .A2(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3148_ (.A1(_1926_),
    .A2(_0290_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3149_ (.A1(_1934_),
    .A2(_0291_),
    .B(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3150_ (.A1(_0289_),
    .A2(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3151_ (.A1(_0289_),
    .A2(_0293_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3152_ (.A1(_0288_),
    .A2(_0294_),
    .B(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3153_ (.A1(_0266_),
    .A2(_0267_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3154_ (.I(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3155_ (.A1(_0274_),
    .A2(_0275_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3156_ (.I(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3157_ (.A1(_0277_),
    .A2(_0296_),
    .B(_0298_),
    .C(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3158_ (.I(_0251_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3159_ (.A1(_0302_),
    .A2(_0258_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3160_ (.I(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3161_ (.A1(_0261_),
    .A2(_0269_),
    .A3(_0301_),
    .A4(_0304_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3162_ (.A1(_0237_),
    .A2(_0243_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3163_ (.I(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3164_ (.A1(_0260_),
    .A2(_0305_),
    .B(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3165_ (.A1(_0230_),
    .A2(_0234_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3166_ (.I(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3167_ (.A1(_0244_),
    .A2(_0308_),
    .B(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3168_ (.A1(_0223_),
    .A2(_0228_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3169_ (.A1(_0236_),
    .A2(_0311_),
    .B(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3170_ (.A1(_0214_),
    .A2(_0219_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3171_ (.I(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3172_ (.A1(_0229_),
    .A2(_0313_),
    .B(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3173_ (.I(_2037_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3174_ (.I(\Control_Unit.T[12] ),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3175_ (.I(_2041_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3176_ (.I(_0319_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3177_ (.A1(_0317_),
    .A2(_0318_),
    .A3(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3178_ (.I(_1713_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3179_ (.A1(_0222_),
    .A2(_0213_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3180_ (.A1(_0222_),
    .A2(_0213_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3181_ (.A1(_0322_),
    .A2(_0323_),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3182_ (.A1(_0321_),
    .A2(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3183_ (.A1(_0221_),
    .A2(_0316_),
    .A3(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3184_ (.I(_0229_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3185_ (.I(_0244_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3186_ (.A1(_0261_),
    .A2(_0269_),
    .A3(_0301_),
    .A4(_0304_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3187_ (.A1(_0259_),
    .A2(_0330_),
    .B(_0306_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3188_ (.A1(_0329_),
    .A2(_0331_),
    .B(_0309_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3189_ (.I(_0312_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3190_ (.A1(_0235_),
    .A2(_0332_),
    .B(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3191_ (.A1(_0328_),
    .A2(_0334_),
    .B(_0314_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3192_ (.I(_0326_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3193_ (.A1(_0220_),
    .A2(_0335_),
    .B(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3194_ (.I(\Control_Unit.Rc ),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3195_ (.A1(_0338_),
    .A2(\Control_Unit.Mt ),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3196_ (.I(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3197_ (.I(_0340_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3198_ (.I(\Control_Unit.Mt ),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3199_ (.I(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3200_ (.I(_0343_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3201_ (.I(\Control_Unit.T[12] ),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3202_ (.A1(_0327_),
    .A2(_0337_),
    .A3(_0341_),
    .B1(_0344_),
    .B2(_0345_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3203_ (.I(_0339_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3204_ (.I(_0346_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3205_ (.A1(_0321_),
    .A2(_0325_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3206_ (.I(\Control_Unit.T[13] ),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3207_ (.A1(_0319_),
    .A2(_0349_),
    .A3(_1881_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3208_ (.I(_1711_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3209_ (.A1(_0317_),
    .A2(_0318_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3210_ (.A1(_0317_),
    .A2(_0318_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3211_ (.A1(_0351_),
    .A2(_0352_),
    .B(_0353_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3212_ (.A1(_0350_),
    .A2(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3213_ (.A1(_0348_),
    .A2(_0337_),
    .A3(_0355_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3214_ (.A1(_0321_),
    .A2(_0325_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3215_ (.A1(_0221_),
    .A2(_0316_),
    .B(_0326_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3216_ (.I(_0355_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3217_ (.A1(_0357_),
    .A2(_0358_),
    .B(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3218_ (.I(\Control_Unit.T[13] ),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3219_ (.A1(_0347_),
    .A2(_0356_),
    .A3(_0360_),
    .B1(_0344_),
    .B2(_0361_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3220_ (.I(\Control_Unit.T[14] ),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3221_ (.I(_0343_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3222_ (.A1(_0350_),
    .A2(_0354_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3223_ (.A1(_0348_),
    .A2(_0337_),
    .B(_0355_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3224_ (.I(\Control_Unit.T[14] ),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3225_ (.A1(_1881_),
    .A2(_0366_),
    .A3(_2177_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3226_ (.A1(_0320_),
    .A2(_0349_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3227_ (.A1(_0320_),
    .A2(_0349_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3228_ (.A1(_1889_),
    .A2(_0368_),
    .B(_0369_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3229_ (.A1(_0367_),
    .A2(_0370_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3230_ (.I(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3231_ (.A1(_0364_),
    .A2(_0365_),
    .B(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3232_ (.I(_0364_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3233_ (.I(\Control_Unit.Mt ),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3234_ (.A1(\Control_Unit.Rc ),
    .A2(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3235_ (.I(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3236_ (.I(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3237_ (.A1(_0374_),
    .A2(_0360_),
    .A3(_0371_),
    .B(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3238_ (.A1(_0362_),
    .A2(_0363_),
    .B1(_0373_),
    .B2(_0379_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3239_ (.I(_0346_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3240_ (.A1(_0367_),
    .A2(_0370_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3241_ (.I(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3242_ (.I(_1707_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3243_ (.I(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3244_ (.I(\Control_Unit.T[15] ),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3245_ (.A1(_2176_),
    .A2(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3246_ (.A1(_0384_),
    .A2(_0386_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3247_ (.I(_1710_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3248_ (.A1(_1882_),
    .A2(_0366_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3249_ (.A1(_1882_),
    .A2(_0366_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3250_ (.A1(_0388_),
    .A2(_0389_),
    .B(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3251_ (.A1(_0387_),
    .A2(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3252_ (.A1(_0382_),
    .A2(_0373_),
    .A3(_0392_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3253_ (.A1(_0374_),
    .A2(_0360_),
    .B(_0371_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3254_ (.I(_0392_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3255_ (.A1(_0381_),
    .A2(_0394_),
    .B(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3256_ (.I(_0343_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3257_ (.I(_0385_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3258_ (.A1(_0380_),
    .A2(_0393_),
    .A3(_0396_),
    .B1(_0397_),
    .B2(_0398_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3259_ (.I(\Control_Unit.T[16] ),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3260_ (.A1(_0387_),
    .A2(_0391_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3261_ (.A1(_0382_),
    .A2(_0373_),
    .B(_0392_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3262_ (.A1(_0400_),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3263_ (.I(\Control_Unit.T[16] ),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3264_ (.A1(_0384_),
    .A2(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3265_ (.A1(_0384_),
    .A2(_0403_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3266_ (.A1(_0404_),
    .A2(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3267_ (.A1(_1966_),
    .A2(_0386_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3268_ (.A1(_0388_),
    .A2(_0398_),
    .B(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3269_ (.A1(_0406_),
    .A2(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3270_ (.I(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3271_ (.A1(_0402_),
    .A2(_0410_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3272_ (.A1(_0402_),
    .A2(_0410_),
    .B(_0378_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3273_ (.A1(_0399_),
    .A2(_0363_),
    .B1(_0411_),
    .B2(_0412_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3274_ (.I(\Control_Unit.T[17] ),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3275_ (.I(_0404_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3276_ (.A1(_0414_),
    .A2(_0405_),
    .A3(_0408_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3277_ (.A1(_0387_),
    .A2(_0391_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3278_ (.A1(_0416_),
    .A2(_0396_),
    .B(_0410_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3279_ (.A1(_0415_),
    .A2(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3280_ (.A1(_0413_),
    .A2(_0414_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3281_ (.A1(_0418_),
    .A2(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3282_ (.A1(_0413_),
    .A2(_0363_),
    .B1(_0341_),
    .B2(_0420_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3283_ (.I(\Control_Unit.Rc ),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3284_ (.I(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3285_ (.A1(_0414_),
    .A2(_0415_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3286_ (.A1(\Control_Unit.T[17] ),
    .A2(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3287_ (.A1(_0409_),
    .A2(_0419_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3288_ (.A1(_0416_),
    .A2(_0396_),
    .B(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3289_ (.I(\Control_Unit.T[18] ),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3290_ (.A1(_0424_),
    .A2(_0426_),
    .B(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3291_ (.A1(_0422_),
    .A2(_0428_),
    .B(_0342_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3292_ (.I(\Control_Unit.T[18] ),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3293_ (.A1(_0424_),
    .A2(_0426_),
    .B(_0346_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3294_ (.A1(_0430_),
    .A2(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3295_ (.A1(_0429_),
    .A2(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3296_ (.I(_0433_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3297_ (.A1(_0424_),
    .A2(_0426_),
    .B(_0427_),
    .C(_0346_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3298_ (.I(\Control_Unit.T[19] ),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3299_ (.I0(_0434_),
    .I1(_0429_),
    .S(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3300_ (.I(_0436_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3301_ (.A1(_0430_),
    .A2(_0435_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3302_ (.I(\Control_Unit.T[20] ),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3303_ (.A1(_0424_),
    .A2(_0426_),
    .B(_0437_),
    .C(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3304_ (.A1(_0380_),
    .A2(_0439_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3305_ (.A1(_0435_),
    .A2(_0434_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3306_ (.A1(_0344_),
    .A2(_0440_),
    .B1(_0441_),
    .B2(_0438_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3307_ (.I(_0376_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3308_ (.A1(_0442_),
    .A2(_0439_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3309_ (.A1(_0422_),
    .A2(_0439_),
    .B(_0343_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3310_ (.I(\Control_Unit.T[21] ),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3311_ (.I0(_0443_),
    .I1(_0444_),
    .S(_0445_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3312_ (.I(_0446_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3313_ (.I(\Control_Unit.T[22] ),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3314_ (.A1(_0414_),
    .A2(_0415_),
    .B(_0413_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3315_ (.A1(_0410_),
    .A2(_0419_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3316_ (.A1(_0400_),
    .A2(_0401_),
    .B(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3317_ (.A1(_0430_),
    .A2(_0435_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3318_ (.A1(\Control_Unit.T[20] ),
    .A2(_0445_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3319_ (.A1(_0448_),
    .A2(_0450_),
    .B(_0451_),
    .C(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3320_ (.A1(_0447_),
    .A2(_0453_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3321_ (.A1(_0447_),
    .A2(_0453_),
    .B(_0442_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3322_ (.A1(_0447_),
    .A2(_0344_),
    .B1(_0454_),
    .B2(_0455_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3323_ (.I(\Control_Unit.T[23] ),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3324_ (.I(\Control_Unit.T[22] ),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3325_ (.A1(_0445_),
    .A2(_0457_),
    .A3(_0378_),
    .A4(_0439_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3326_ (.I(_0375_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3327_ (.A1(_0456_),
    .A2(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3328_ (.A1(_0456_),
    .A2(_0458_),
    .B1(_0460_),
    .B2(_0455_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3329_ (.A1(_0457_),
    .A2(\Control_Unit.T[23] ),
    .A3(_0451_),
    .A4(_0452_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3330_ (.A1(_0416_),
    .A2(_0396_),
    .B(_0425_),
    .C(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3331_ (.A1(_0448_),
    .A2(_0461_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3332_ (.I(\Control_Unit.T[24] ),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3333_ (.A1(_0462_),
    .A2(_0463_),
    .B(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3334_ (.A1(_0422_),
    .A2(_0465_),
    .B(_0342_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3335_ (.A1(_0425_),
    .A2(_0461_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3336_ (.A1(_0400_),
    .A2(_0401_),
    .B(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3337_ (.I(_0463_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3338_ (.A1(_0468_),
    .A2(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3339_ (.A1(_0380_),
    .A2(_0470_),
    .B(_0464_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3340_ (.A1(_0466_),
    .A2(_0471_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3341_ (.I(_0472_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3342_ (.A1(_0377_),
    .A2(_0465_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3343_ (.I(\Control_Unit.T[25] ),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3344_ (.I0(_0473_),
    .I1(_0466_),
    .S(_0474_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3345_ (.I(_0475_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3346_ (.A1(\Control_Unit.T[24] ),
    .A2(_0474_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3347_ (.I(\Control_Unit.T[26] ),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3348_ (.I(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3349_ (.A1(_0462_),
    .A2(_0463_),
    .B(_0476_),
    .C(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3350_ (.A1(_0422_),
    .A2(_0479_),
    .B(_0342_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3351_ (.A1(_0380_),
    .A2(_0470_),
    .A3(_0476_),
    .B(_0478_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3352_ (.A1(_0480_),
    .A2(_0481_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3353_ (.I(_0482_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3354_ (.A1(_0377_),
    .A2(_0479_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3355_ (.I(\Control_Unit.T[27] ),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3356_ (.I0(_0483_),
    .I1(_0480_),
    .S(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3357_ (.I(_0485_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3358_ (.I(\Control_Unit.T[28] ),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3359_ (.A1(_0477_),
    .A2(_0484_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3360_ (.A1(_0462_),
    .A2(_0463_),
    .B(_0476_),
    .C(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3361_ (.A1(_0442_),
    .A2(_0488_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3362_ (.I(_0338_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3363_ (.A1(_0476_),
    .A2(_0487_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3364_ (.I(\Control_Unit.T[28] ),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3365_ (.A1(_0468_),
    .A2(_0469_),
    .B(_0491_),
    .C(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3366_ (.A1(_0490_),
    .A2(_0493_),
    .B(_0459_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3367_ (.A1(_0486_),
    .A2(_0489_),
    .B(_0494_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3368_ (.I(\Control_Unit.T[29] ),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3369_ (.A1(_0492_),
    .A2(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3370_ (.A1(_0495_),
    .A2(_0494_),
    .B1(_0489_),
    .B2(_0496_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3371_ (.I(\Control_Unit.T[30] ),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3372_ (.A1(_0486_),
    .A2(_0495_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3373_ (.A1(_0468_),
    .A2(_0469_),
    .B(_0491_),
    .C(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3374_ (.I(\Control_Unit.T[30] ),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3375_ (.A1(_0500_),
    .A2(_0459_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3376_ (.A1(_0497_),
    .A2(_0499_),
    .B(_0442_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3377_ (.A1(_0497_),
    .A2(_0499_),
    .B1(_0501_),
    .B2(_0502_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3378_ (.I(\Control_Unit.T[31] ),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3379_ (.A1(_0500_),
    .A2(_0378_),
    .A3(_0488_),
    .A4(_0498_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3380_ (.A1(_0503_),
    .A2(_0459_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3381_ (.A1(_0503_),
    .A2(_0504_),
    .B1(_0505_),
    .B2(_0502_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3382_ (.I(_2153_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3383_ (.I(\Control_Unit.Rcont ),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3384_ (.I(_0507_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3385_ (.A1(_0506_),
    .A2(_0508_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3386_ (.A1(_0508_),
    .A2(_2145_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3387_ (.I(_0507_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3388_ (.A1(_0509_),
    .A2(_1816_),
    .A3(_1817_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3389_ (.A1(_0508_),
    .A2(_2265_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3390_ (.A1(_0508_),
    .A2(_2068_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3391_ (.A1(_0509_),
    .A2(_1844_),
    .A3(_1842_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3392_ (.I(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3393_ (.A1(_0510_),
    .A2(_2061_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3394_ (.I(\Control_Unit.Rcont ),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3395_ (.A1(_0511_),
    .A2(_2118_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3396_ (.I(_0512_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3397_ (.A1(_0510_),
    .A2(_1758_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3398_ (.A1(_0510_),
    .A2(_1864_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3399_ (.A1(_0510_),
    .A2(_1863_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3400_ (.A1(_0509_),
    .A2(_2191_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3401_ (.A1(_0511_),
    .A2(_1877_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3402_ (.I(_0513_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3403_ (.A1(_0511_),
    .A2(_2173_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3404_ (.I(_0514_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3405_ (.A1(_0511_),
    .A2(_2174_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3406_ (.I(_0515_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3407_ (.A1(\Control_Unit.Rcont ),
    .A2(_1730_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3408_ (.I(_0516_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3409_ (.I(net19),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3410_ (.I(\Control_Unit.Mx ),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3411_ (.I(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3412_ (.I(\Control_Unit.Rx ),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3413_ (.A1(_0520_),
    .A2(\Control_Unit.Mx ),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3414_ (.I(_0521_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3415_ (.I(_0522_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3416_ (.I(_0523_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3417_ (.I(_2014_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3418_ (.A1(\Control_Unit.Q[0] ),
    .A2(\Control_Unit.T[0] ),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3419_ (.A1(_0525_),
    .A2(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3420_ (.A1(_0517_),
    .A2(_0519_),
    .B1(_0524_),
    .B2(_0527_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3421_ (.I(\Control_Unit.Mx ),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3422_ (.I(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3423_ (.I(net30),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3424_ (.I(\Control_Unit.Q[0] ),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3425_ (.I(_0278_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3426_ (.I(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3427_ (.A1(_0531_),
    .A2(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3428_ (.A1(_2014_),
    .A2(_0526_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3429_ (.I(\Control_Unit.T[1] ),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3430_ (.A1(\Control_Unit.C[1] ),
    .A2(\Control_Unit.Q[1] ),
    .A3(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3431_ (.A1(_0534_),
    .A2(_0535_),
    .A3(_0537_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3432_ (.A1(_0529_),
    .A2(_0530_),
    .B1(_0524_),
    .B2(_0538_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3433_ (.I(_0521_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3434_ (.I(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3435_ (.I(\Control_Unit.C[2] ),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3436_ (.I(\Control_Unit.Q[2] ),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3437_ (.A1(_0541_),
    .A2(_0542_),
    .A3(\Control_Unit.T[2] ),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3438_ (.I(\Control_Unit.Q[1] ),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3439_ (.A1(_2013_),
    .A2(_0536_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3440_ (.A1(_2013_),
    .A2(_0536_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3441_ (.A1(_0544_),
    .A2(_0545_),
    .B(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3442_ (.A1(_0543_),
    .A2(_0547_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3443_ (.I(_0531_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3444_ (.A1(_0549_),
    .A2(_0278_),
    .A3(_0537_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3445_ (.A1(_0549_),
    .A2(_0278_),
    .B(_0537_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3446_ (.A1(_0535_),
    .A2(_0550_),
    .B(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3447_ (.A1(_0548_),
    .A2(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3448_ (.A1(_0548_),
    .A2(_0552_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3449_ (.I(net41),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3450_ (.A1(_0540_),
    .A2(_0553_),
    .A3(_0554_),
    .B1(_0555_),
    .B2(_0519_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3451_ (.A1(_2016_),
    .A2(\Control_Unit.T[2] ),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3452_ (.I(\Control_Unit.Q[3] ),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3453_ (.A1(\Control_Unit.C[3] ),
    .A2(\Control_Unit.T[3] ),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3454_ (.A1(_0557_),
    .A2(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3455_ (.A1(_2016_),
    .A2(_0290_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3456_ (.A1(_0542_),
    .A2(_0556_),
    .B(_0559_),
    .C(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3457_ (.A1(_0542_),
    .A2(_0556_),
    .B(_0560_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3458_ (.I(_0557_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3459_ (.A1(_0563_),
    .A2(_0558_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3460_ (.A1(_0563_),
    .A2(_0558_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3461_ (.A1(_0562_),
    .A2(_0564_),
    .A3(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3462_ (.A1(_0543_),
    .A2(_0547_),
    .B1(_0561_),
    .B2(_0566_),
    .C(_0553_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3463_ (.A1(_0543_),
    .A2(_0547_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3464_ (.A1(_0548_),
    .A2(_0552_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3465_ (.I(_0561_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3466_ (.A1(_0562_),
    .A2(_0564_),
    .A3(_0565_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3467_ (.A1(_0568_),
    .A2(_0569_),
    .B(_0570_),
    .C(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3468_ (.I(net44),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3469_ (.A1(_0540_),
    .A2(_0567_),
    .A3(_0572_),
    .B1(_0573_),
    .B2(_0519_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3470_ (.I(net45),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3471_ (.A1(\Control_Unit.T[4] ),
    .A2(_2008_),
    .A3(\Control_Unit.Q[4] ),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3472_ (.A1(_2015_),
    .A2(_0270_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3473_ (.A1(_0563_),
    .A2(_0558_),
    .B(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3474_ (.A1(_0575_),
    .A2(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3475_ (.A1(_0543_),
    .A2(_0547_),
    .B1(_0548_),
    .B2(_0552_),
    .C(_0571_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3476_ (.A1(_0570_),
    .A2(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3477_ (.A1(_0578_),
    .A2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3478_ (.A1(_0529_),
    .A2(_0574_),
    .B1(_0524_),
    .B2(_0581_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3479_ (.I(_0518_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3480_ (.I(net46),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3481_ (.I(\Control_Unit.Q[5] ),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3482_ (.A1(\Control_Unit.T[5] ),
    .A2(_2006_),
    .A3(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3483_ (.I(\Control_Unit.Q[4] ),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3484_ (.A1(_0262_),
    .A2(_2009_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3485_ (.A1(_0262_),
    .A2(_2009_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3486_ (.A1(_0586_),
    .A2(_0587_),
    .B(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3487_ (.A1(_0585_),
    .A2(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3488_ (.A1(_0585_),
    .A2(_0589_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3489_ (.A1(_0590_),
    .A2(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3490_ (.A1(_0576_),
    .A2(_0564_),
    .B(_0575_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3491_ (.A1(_0578_),
    .A2(_0580_),
    .B(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3492_ (.A1(_0592_),
    .A2(_0594_),
    .B(_0539_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3493_ (.A1(_0592_),
    .A2(_0594_),
    .B(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3494_ (.A1(_0582_),
    .A2(_0583_),
    .B(_0596_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3495_ (.I(net47),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3496_ (.I(\Control_Unit.T[6] ),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3497_ (.I(\Control_Unit.Q[6] ),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3498_ (.A1(_0598_),
    .A2(\Control_Unit.C[6] ),
    .A3(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3499_ (.A1(_0254_),
    .A2(_2007_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3500_ (.A1(_0254_),
    .A2(_2007_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3501_ (.A1(_0584_),
    .A2(_0601_),
    .B(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3502_ (.A1(_0600_),
    .A2(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3503_ (.A1(_0578_),
    .A2(_0590_),
    .A3(_0591_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3504_ (.A1(_0585_),
    .A2(_0589_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3505_ (.A1(_0593_),
    .A2(_0606_),
    .B(_0591_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3506_ (.A1(_0570_),
    .A2(_0579_),
    .A3(_0605_),
    .B(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3507_ (.A1(_0604_),
    .A2(_0608_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3508_ (.A1(_0529_),
    .A2(_0597_),
    .B1(_0524_),
    .B2(_0609_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3509_ (.I(net48),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3510_ (.I(\Control_Unit.Q[7] ),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3511_ (.A1(\Control_Unit.T[7] ),
    .A2(\Control_Unit.C[7] ),
    .A3(_0611_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3512_ (.I(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3513_ (.A1(_0246_),
    .A2(_2011_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3514_ (.A1(_0246_),
    .A2(_2011_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3515_ (.A1(_0599_),
    .A2(_0614_),
    .B(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3516_ (.A1(_0613_),
    .A2(_0616_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3517_ (.A1(_0600_),
    .A2(_0603_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3518_ (.A1(_0604_),
    .A2(_0608_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3519_ (.A1(_0618_),
    .A2(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3520_ (.A1(_0617_),
    .A2(_0620_),
    .B(_0539_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3521_ (.A1(_0617_),
    .A2(_0620_),
    .B(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3522_ (.A1(_0582_),
    .A2(_0610_),
    .B(_0622_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3523_ (.I(_0528_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3524_ (.I(net49),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3525_ (.I(_0523_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3526_ (.A1(_0604_),
    .A2(_0617_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3527_ (.A1(_0570_),
    .A2(_0579_),
    .A3(_0605_),
    .A4(_0626_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3528_ (.A1(_0613_),
    .A2(_0616_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3529_ (.A1(_0613_),
    .A2(_0616_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3530_ (.A1(_0618_),
    .A2(_0628_),
    .B1(_0626_),
    .B2(_0607_),
    .C(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3531_ (.A1(_0627_),
    .A2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3532_ (.A1(\Control_Unit.T[8] ),
    .A2(_2001_),
    .A3(\Control_Unit.Q[8] ),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3533_ (.A1(\Control_Unit.T[7] ),
    .A2(_2010_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3534_ (.A1(_0240_),
    .A2(_2010_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3535_ (.A1(_0611_),
    .A2(_0633_),
    .B(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3536_ (.A1(_0632_),
    .A2(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3537_ (.I(_0636_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3538_ (.A1(_0631_),
    .A2(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3539_ (.A1(_0623_),
    .A2(_0624_),
    .B1(_0625_),
    .B2(_0638_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3540_ (.I(net50),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3541_ (.A1(\Control_Unit.T[9] ),
    .A2(_2000_),
    .A3(\Control_Unit.Q[9] ),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3542_ (.A1(\Control_Unit.T[8] ),
    .A2(\Control_Unit.C[8] ),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3543_ (.A1(_0231_),
    .A2(\Control_Unit.C[8] ),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3544_ (.A1(\Control_Unit.Q[8] ),
    .A2(_0641_),
    .B(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3545_ (.A1(_0640_),
    .A2(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3546_ (.A1(_0632_),
    .A2(_0635_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3547_ (.A1(_0631_),
    .A2(_0636_),
    .B(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3548_ (.A1(_0644_),
    .A2(_0646_),
    .B(_0539_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3549_ (.A1(_0644_),
    .A2(_0646_),
    .B(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3550_ (.A1(_0582_),
    .A2(_0639_),
    .B(_0648_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3551_ (.I(net20),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3552_ (.A1(_0627_),
    .A2(_0630_),
    .B(_0637_),
    .C(_0644_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3553_ (.A1(_0640_),
    .A2(_0643_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3554_ (.A1(_0640_),
    .A2(_0643_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3555_ (.A1(_0645_),
    .A2(_0651_),
    .B(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3556_ (.I(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3557_ (.A1(_0650_),
    .A2(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3558_ (.A1(\Control_Unit.T[10] ),
    .A2(_2004_),
    .A3(\Control_Unit.Q[10] ),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3559_ (.A1(\Control_Unit.T[9] ),
    .A2(\Control_Unit.C[9] ),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3560_ (.A1(_0225_),
    .A2(\Control_Unit.C[9] ),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3561_ (.A1(\Control_Unit.Q[9] ),
    .A2(_0657_),
    .B(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3562_ (.A1(_0656_),
    .A2(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3563_ (.A1(_0655_),
    .A2(_0660_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3564_ (.A1(_0623_),
    .A2(_0649_),
    .B1(_0625_),
    .B2(_0661_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3565_ (.I(_0518_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3566_ (.I(net21),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3567_ (.A1(\Control_Unit.T[11] ),
    .A2(_2002_),
    .A3(\Control_Unit.Q[11] ),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3568_ (.A1(\Control_Unit.T[10] ),
    .A2(\Control_Unit.C[10] ),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3569_ (.A1(\Control_Unit.T[10] ),
    .A2(\Control_Unit.C[10] ),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3570_ (.A1(\Control_Unit.Q[10] ),
    .A2(_0665_),
    .B(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3571_ (.A1(_0664_),
    .A2(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3572_ (.I(_0660_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3573_ (.A1(_0656_),
    .A2(_0659_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3574_ (.A1(_0655_),
    .A2(_0669_),
    .B(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3575_ (.I(_0522_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3576_ (.A1(_0668_),
    .A2(_0671_),
    .B(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3577_ (.A1(_0668_),
    .A2(_0671_),
    .B(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3578_ (.A1(_0662_),
    .A2(_0663_),
    .B(_0674_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3579_ (.I(net22),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3580_ (.A1(_0650_),
    .A2(_0654_),
    .B(_0660_),
    .C(_0668_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3581_ (.I(_0667_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3582_ (.A1(_0664_),
    .A2(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3583_ (.A1(_0664_),
    .A2(_0677_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3584_ (.A1(_0670_),
    .A2(_0678_),
    .B(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3585_ (.I(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3586_ (.A1(_0676_),
    .A2(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3587_ (.A1(_0345_),
    .A2(\Control_Unit.C[12] ),
    .A3(\Control_Unit.Q[12] ),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3588_ (.A1(\Control_Unit.T[11] ),
    .A2(_2002_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3589_ (.A1(\Control_Unit.T[11] ),
    .A2(_2002_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3590_ (.A1(\Control_Unit.Q[11] ),
    .A2(_0684_),
    .B(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3591_ (.A1(_0683_),
    .A2(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3592_ (.I(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3593_ (.A1(_0682_),
    .A2(_0688_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3594_ (.A1(_0623_),
    .A2(_0675_),
    .B1(_0625_),
    .B2(_0689_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3595_ (.I(net23),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3596_ (.A1(_0361_),
    .A2(\Control_Unit.C[13] ),
    .A3(\Control_Unit.Q[13] ),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3597_ (.A1(\Control_Unit.T[12] ),
    .A2(_2019_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3598_ (.A1(_0318_),
    .A2(_2019_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3599_ (.A1(\Control_Unit.Q[12] ),
    .A2(_0692_),
    .B(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3600_ (.A1(_0691_),
    .A2(_0694_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3601_ (.A1(_0683_),
    .A2(_0686_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3602_ (.A1(_0682_),
    .A2(_0687_),
    .B(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3603_ (.A1(_0695_),
    .A2(_0697_),
    .B(_0672_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3604_ (.A1(_0695_),
    .A2(_0697_),
    .B(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3605_ (.A1(_0662_),
    .A2(_0690_),
    .B(_0699_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3606_ (.I(net24),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3607_ (.A1(_0676_),
    .A2(_0681_),
    .B(_0688_),
    .C(_0695_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3608_ (.A1(_0691_),
    .A2(_0694_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3609_ (.A1(_0691_),
    .A2(_0694_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3610_ (.A1(_0696_),
    .A2(_0702_),
    .B(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3611_ (.I(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3612_ (.A1(_0701_),
    .A2(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3613_ (.A1(_0362_),
    .A2(\Control_Unit.C[14] ),
    .A3(\Control_Unit.Q[14] ),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3614_ (.A1(\Control_Unit.T[13] ),
    .A2(_2018_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3615_ (.A1(_0349_),
    .A2(_2018_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3616_ (.A1(\Control_Unit.Q[13] ),
    .A2(_0708_),
    .B(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3617_ (.A1(_0707_),
    .A2(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3618_ (.A1(_0706_),
    .A2(_0711_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3619_ (.A1(_0623_),
    .A2(_0700_),
    .B1(_0625_),
    .B2(_0712_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3620_ (.I(net25),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3621_ (.I(\Control_Unit.Q[15] ),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3622_ (.A1(\Control_Unit.T[15] ),
    .A2(\Control_Unit.C[15] ),
    .A3(_0714_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3623_ (.A1(\Control_Unit.T[14] ),
    .A2(_2021_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3624_ (.A1(_0366_),
    .A2(_2021_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3625_ (.A1(\Control_Unit.Q[14] ),
    .A2(_0716_),
    .B(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3626_ (.A1(_0715_),
    .A2(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3627_ (.I(_0711_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3628_ (.A1(_0707_),
    .A2(_0710_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3629_ (.A1(_0706_),
    .A2(_0720_),
    .B(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3630_ (.A1(_0719_),
    .A2(_0722_),
    .B(_0672_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3631_ (.A1(_0719_),
    .A2(_0722_),
    .B(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3632_ (.A1(_0662_),
    .A2(_0713_),
    .B(_0724_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3633_ (.I(_0528_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3634_ (.I(net26),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3635_ (.I(_0523_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3636_ (.A1(_0701_),
    .A2(_0705_),
    .B(_0711_),
    .C(_0719_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3637_ (.I(_0718_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3638_ (.A1(_0715_),
    .A2(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3639_ (.A1(_0715_),
    .A2(_0729_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3640_ (.A1(_0721_),
    .A2(_0730_),
    .B(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3641_ (.I(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3642_ (.A1(_0728_),
    .A2(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3643_ (.A1(_0399_),
    .A2(\Control_Unit.C[16] ),
    .A3(\Control_Unit.Q[16] ),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3644_ (.A1(_0385_),
    .A2(_2020_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3645_ (.A1(_0385_),
    .A2(_2020_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3646_ (.A1(_0714_),
    .A2(_0736_),
    .B(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3647_ (.A1(_0735_),
    .A2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3648_ (.I(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3649_ (.A1(_0734_),
    .A2(_0740_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3650_ (.A1(_0725_),
    .A2(_0726_),
    .B1(_0727_),
    .B2(_0741_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3651_ (.I(net27),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3652_ (.I(\Control_Unit.Q[17] ),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3653_ (.A1(_0413_),
    .A2(\Control_Unit.C[17] ),
    .A3(_0743_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3654_ (.A1(_0403_),
    .A2(\Control_Unit.C[16] ),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3655_ (.A1(_0403_),
    .A2(_1989_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3656_ (.A1(\Control_Unit.Q[16] ),
    .A2(_0745_),
    .B(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3657_ (.A1(_0744_),
    .A2(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3658_ (.A1(_0735_),
    .A2(_0738_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3659_ (.A1(_0734_),
    .A2(_0739_),
    .B(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3660_ (.A1(_0748_),
    .A2(_0750_),
    .B(_0672_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3661_ (.A1(_0748_),
    .A2(_0750_),
    .B(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3662_ (.A1(_0662_),
    .A2(_0742_),
    .B(_0752_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3663_ (.I(net28),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3664_ (.A1(_0728_),
    .A2(_0733_),
    .B(_0740_),
    .C(_0748_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3665_ (.A1(_0744_),
    .A2(_0747_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3666_ (.A1(_0749_),
    .A2(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3667_ (.A1(_0744_),
    .A2(_0747_),
    .B(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3668_ (.A1(_0754_),
    .A2(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3669_ (.A1(_0427_),
    .A2(\Control_Unit.C[18] ),
    .A3(\Control_Unit.Q[18] ),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3670_ (.A1(\Control_Unit.T[17] ),
    .A2(_1987_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3671_ (.A1(\Control_Unit.T[17] ),
    .A2(_1987_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3672_ (.A1(_0743_),
    .A2(_0760_),
    .B(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3673_ (.A1(_0759_),
    .A2(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3674_ (.A1(_0758_),
    .A2(_0763_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3675_ (.A1(_0725_),
    .A2(_0753_),
    .B1(_0727_),
    .B2(_0764_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3676_ (.I(_0518_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3677_ (.I(net29),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3678_ (.A1(\Control_Unit.T[19] ),
    .A2(\Control_Unit.C[19] ),
    .A3(\Control_Unit.Q[19] ),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3679_ (.I(\Control_Unit.Q[18] ),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3680_ (.A1(\Control_Unit.T[18] ),
    .A2(_1992_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3681_ (.A1(_0430_),
    .A2(_1992_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3682_ (.A1(_0768_),
    .A2(_0769_),
    .B(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3683_ (.A1(_0767_),
    .A2(_0771_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3684_ (.A1(_0759_),
    .A2(_0762_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3685_ (.A1(_0754_),
    .A2(_0757_),
    .B(_0763_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3686_ (.A1(_0773_),
    .A2(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3687_ (.I(_0522_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3688_ (.A1(_0772_),
    .A2(_0775_),
    .B(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3689_ (.A1(_0772_),
    .A2(_0775_),
    .B(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3690_ (.A1(_0765_),
    .A2(_0766_),
    .B(_0778_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3691_ (.I(net31),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3692_ (.A1(_0754_),
    .A2(_0757_),
    .B(_0763_),
    .C(_0772_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3693_ (.I(_0771_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3694_ (.A1(_0767_),
    .A2(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3695_ (.A1(_0767_),
    .A2(_0781_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3696_ (.A1(_0773_),
    .A2(_0782_),
    .B(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3697_ (.I(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3698_ (.A1(_0780_),
    .A2(_0785_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3699_ (.A1(_0438_),
    .A2(\Control_Unit.C[20] ),
    .A3(\Control_Unit.Q[20] ),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3700_ (.I(\Control_Unit.Q[19] ),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3701_ (.A1(\Control_Unit.T[19] ),
    .A2(_1990_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3702_ (.A1(\Control_Unit.T[19] ),
    .A2(_1990_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3703_ (.A1(_0788_),
    .A2(_0789_),
    .B(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3704_ (.A1(_0787_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3705_ (.I(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3706_ (.A1(_0786_),
    .A2(_0793_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3707_ (.A1(_0725_),
    .A2(_0779_),
    .B1(_0727_),
    .B2(_0794_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3708_ (.I(net32),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3709_ (.A1(\Control_Unit.T[21] ),
    .A2(\Control_Unit.C[21] ),
    .A3(\Control_Unit.Q[21] ),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3710_ (.I(\Control_Unit.Q[20] ),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3711_ (.A1(\Control_Unit.T[20] ),
    .A2(\Control_Unit.C[20] ),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3712_ (.A1(\Control_Unit.T[20] ),
    .A2(_1983_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3713_ (.A1(_0797_),
    .A2(_0798_),
    .B(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3714_ (.A1(_0796_),
    .A2(_0800_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3715_ (.A1(_0787_),
    .A2(_0791_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3716_ (.A1(_0786_),
    .A2(_0792_),
    .B(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3717_ (.A1(_0801_),
    .A2(_0803_),
    .B(_0776_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3718_ (.A1(_0801_),
    .A2(_0803_),
    .B(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3719_ (.A1(_0765_),
    .A2(_0795_),
    .B(_0805_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3720_ (.I(net33),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3721_ (.A1(_0780_),
    .A2(_0785_),
    .B(_0793_),
    .C(_0801_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3722_ (.A1(_0796_),
    .A2(_0800_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3723_ (.A1(_0796_),
    .A2(_0800_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3724_ (.A1(_0802_),
    .A2(_0808_),
    .B(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3725_ (.I(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3726_ (.A1(_0807_),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3727_ (.A1(_0447_),
    .A2(\Control_Unit.C[22] ),
    .A3(\Control_Unit.Q[22] ),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3728_ (.I(\Control_Unit.Q[21] ),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3729_ (.A1(\Control_Unit.T[21] ),
    .A2(_1981_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3730_ (.A1(_0445_),
    .A2(_1981_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3731_ (.A1(_0814_),
    .A2(_0815_),
    .B(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3732_ (.A1(_0813_),
    .A2(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3733_ (.A1(_0812_),
    .A2(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3734_ (.A1(_0725_),
    .A2(_0806_),
    .B1(_0727_),
    .B2(_0819_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3735_ (.I(net34),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3736_ (.A1(_0456_),
    .A2(\Control_Unit.C[23] ),
    .A3(\Control_Unit.Q[23] ),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3737_ (.I(\Control_Unit.Q[22] ),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3738_ (.A1(_0457_),
    .A2(\Control_Unit.C[22] ),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3739_ (.A1(_0457_),
    .A2(\Control_Unit.C[22] ),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3740_ (.A1(_0822_),
    .A2(_0823_),
    .B(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3741_ (.A1(_0821_),
    .A2(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3742_ (.I(_0818_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3743_ (.A1(_0813_),
    .A2(_0817_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3744_ (.A1(_0812_),
    .A2(_0827_),
    .B(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3745_ (.A1(_0826_),
    .A2(_0829_),
    .B(_0776_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3746_ (.A1(_0826_),
    .A2(_0829_),
    .B(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3747_ (.A1(_0765_),
    .A2(_0820_),
    .B(_0831_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3748_ (.I(_0528_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3749_ (.I(net35),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3750_ (.I(_0523_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3751_ (.A1(_0807_),
    .A2(_0811_),
    .B(_0818_),
    .C(_0826_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3752_ (.A1(_0821_),
    .A2(_0825_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3753_ (.A1(_0821_),
    .A2(_0825_),
    .B(_0828_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3754_ (.A1(_0836_),
    .A2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3755_ (.A1(_0835_),
    .A2(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3756_ (.A1(_0464_),
    .A2(\Control_Unit.C[24] ),
    .A3(\Control_Unit.Q[24] ),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3757_ (.I(\Control_Unit.Q[23] ),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3758_ (.A1(\Control_Unit.T[23] ),
    .A2(_1984_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3759_ (.A1(\Control_Unit.T[23] ),
    .A2(_1984_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3760_ (.A1(_0841_),
    .A2(_0842_),
    .B(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3761_ (.A1(_0840_),
    .A2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3762_ (.I(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3763_ (.A1(_0839_),
    .A2(_0846_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3764_ (.A1(_0832_),
    .A2(_0833_),
    .B1(_0834_),
    .B2(_0847_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3765_ (.I(net36),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3766_ (.A1(\Control_Unit.T[25] ),
    .A2(\Control_Unit.C[25] ),
    .A3(\Control_Unit.Q[25] ),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3767_ (.I(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3768_ (.A1(\Control_Unit.T[24] ),
    .A2(_1977_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3769_ (.A1(\Control_Unit.T[24] ),
    .A2(_1977_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3770_ (.A1(\Control_Unit.Q[24] ),
    .A2(_0851_),
    .B(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3771_ (.A1(_0850_),
    .A2(_0853_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3772_ (.A1(_0840_),
    .A2(_0844_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3773_ (.A1(_0839_),
    .A2(_0845_),
    .B(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3774_ (.A1(_0854_),
    .A2(_0856_),
    .B(_0776_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3775_ (.A1(_0854_),
    .A2(_0856_),
    .B(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3776_ (.A1(_0765_),
    .A2(_0848_),
    .B(_0858_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3777_ (.I(net37),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3778_ (.A1(\Control_Unit.T[26] ),
    .A2(\Control_Unit.C[26] ),
    .A3(\Control_Unit.Q[26] ),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3779_ (.A1(_0474_),
    .A2(\Control_Unit.C[25] ),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3780_ (.A1(_0474_),
    .A2(_1976_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3781_ (.A1(\Control_Unit.Q[25] ),
    .A2(_0861_),
    .B(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3782_ (.A1(_0860_),
    .A2(_0863_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3783_ (.A1(_0846_),
    .A2(_0854_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3784_ (.A1(_0850_),
    .A2(_0853_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3785_ (.A1(_0855_),
    .A2(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3786_ (.A1(_0850_),
    .A2(_0853_),
    .B(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3787_ (.A1(_0839_),
    .A2(_0865_),
    .B(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3788_ (.A1(_0864_),
    .A2(_0869_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3789_ (.A1(_0832_),
    .A2(_0859_),
    .B1(_0834_),
    .B2(_0870_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3790_ (.I(_0860_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3791_ (.A1(_0871_),
    .A2(_0863_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3792_ (.I(_0864_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3793_ (.A1(_0873_),
    .A2(_0869_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3794_ (.A1(\Control_Unit.T[27] ),
    .A2(\Control_Unit.C[27] ),
    .A3(\Control_Unit.Q[27] ),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3795_ (.I(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3796_ (.A1(_0477_),
    .A2(\Control_Unit.C[26] ),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3797_ (.A1(_0477_),
    .A2(\Control_Unit.C[26] ),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3798_ (.A1(\Control_Unit.Q[26] ),
    .A2(_0877_),
    .B(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3799_ (.A1(_0876_),
    .A2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3800_ (.A1(_0876_),
    .A2(_0879_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3801_ (.A1(_0880_),
    .A2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3802_ (.A1(_0872_),
    .A2(_0874_),
    .B(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3803_ (.A1(_0872_),
    .A2(_0874_),
    .A3(_0882_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3804_ (.I(net38),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3805_ (.A1(_0540_),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(_0519_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3806_ (.I(net39),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3807_ (.A1(_0873_),
    .A2(_0880_),
    .A3(_0881_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3808_ (.A1(_0865_),
    .A2(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3809_ (.A1(_0835_),
    .A2(_0838_),
    .B(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3810_ (.A1(_0871_),
    .A2(_0863_),
    .A3(_0881_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3811_ (.A1(_0868_),
    .A2(_0887_),
    .B(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3812_ (.A1(_0876_),
    .A2(_0879_),
    .B(_0891_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3813_ (.A1(_0889_),
    .A2(_0892_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3814_ (.A1(_0486_),
    .A2(\Control_Unit.C[28] ),
    .A3(\Control_Unit.Q[28] ),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3815_ (.I(\Control_Unit.Q[27] ),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3816_ (.A1(_0484_),
    .A2(\Control_Unit.C[27] ),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3817_ (.A1(_0484_),
    .A2(\Control_Unit.C[27] ),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3818_ (.A1(_0895_),
    .A2(_0896_),
    .B(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3819_ (.A1(_0894_),
    .A2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3820_ (.A1(_0893_),
    .A2(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3821_ (.A1(_0832_),
    .A2(_0886_),
    .B1(_0834_),
    .B2(_0900_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3822_ (.I(net40),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3823_ (.A1(_0495_),
    .A2(\Control_Unit.C[29] ),
    .A3(\Control_Unit.Q[29] ),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3824_ (.A1(_0492_),
    .A2(\Control_Unit.C[28] ),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3825_ (.A1(_0492_),
    .A2(_1996_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3826_ (.A1(\Control_Unit.Q[28] ),
    .A2(_0903_),
    .B(_0904_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3827_ (.A1(_0902_),
    .A2(_0905_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3828_ (.A1(_0894_),
    .A2(_0898_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3829_ (.A1(_0893_),
    .A2(_0899_),
    .B(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3830_ (.A1(_0906_),
    .A2(_0908_),
    .B(_0522_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3831_ (.A1(_0906_),
    .A2(_0908_),
    .B(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3832_ (.A1(_0529_),
    .A2(_0901_),
    .B(_0910_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3833_ (.I(net42),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3834_ (.I(_0906_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3835_ (.A1(_0889_),
    .A2(_0892_),
    .B(_0899_),
    .C(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3836_ (.A1(_0902_),
    .A2(_0905_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3837_ (.A1(_0902_),
    .A2(_0905_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3838_ (.A1(_0907_),
    .A2(_0914_),
    .B(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3839_ (.A1(_0497_),
    .A2(\Control_Unit.C[30] ),
    .A3(\Control_Unit.Q[30] ),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3840_ (.A1(\Control_Unit.T[29] ),
    .A2(_1995_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3841_ (.A1(\Control_Unit.T[29] ),
    .A2(_1995_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3842_ (.A1(\Control_Unit.Q[29] ),
    .A2(_0918_),
    .B(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3843_ (.A1(_0917_),
    .A2(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3844_ (.A1(_0913_),
    .A2(_0916_),
    .A3(_0921_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3845_ (.A1(_0913_),
    .A2(_0916_),
    .B(_0921_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3846_ (.A1(_0922_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3847_ (.A1(_0832_),
    .A2(_0911_),
    .B1(_0834_),
    .B2(_0924_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3848_ (.A1(_0917_),
    .A2(_0920_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3849_ (.A1(_0925_),
    .A2(_0923_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3850_ (.I(\Control_Unit.Q[30] ),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3851_ (.A1(_0500_),
    .A2(\Control_Unit.C[30] ),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3852_ (.A1(_0500_),
    .A2(\Control_Unit.C[30] ),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3853_ (.A1(_0927_),
    .A2(_0928_),
    .B(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3854_ (.A1(_0503_),
    .A2(\Control_Unit.C[31] ),
    .A3(\Control_Unit.Q[31] ),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3855_ (.A1(_0930_),
    .A2(_0931_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3856_ (.A1(_0926_),
    .A2(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3857_ (.A1(_0926_),
    .A2(_0932_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3858_ (.I(net43),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3859_ (.A1(_0540_),
    .A2(_0933_),
    .A3(_0934_),
    .B1(_0935_),
    .B2(_0582_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3860_ (.I(\Control_Unit.Mq ),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3861_ (.I(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3862_ (.A1(_0338_),
    .A2(\Control_Unit.Mq ),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3863_ (.I(_0938_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3864_ (.I(_0939_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3865_ (.I(_2153_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3866_ (.A1(_0941_),
    .A2(_0549_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3867_ (.A1(_0549_),
    .A2(_0937_),
    .B1(_0940_),
    .B2(_0942_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3868_ (.A1(_0282_),
    .A2(_1804_),
    .A3(_0544_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3869_ (.A1(_0506_),
    .A2(_0531_),
    .B(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3870_ (.I(\Control_Unit.Mq ),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3871_ (.A1(\Control_Unit.Rc ),
    .A2(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3872_ (.I(_0946_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3873_ (.A1(_1813_),
    .A2(_0531_),
    .A3(_0943_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3874_ (.A1(_0947_),
    .A2(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3875_ (.I(_0945_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3876_ (.I(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3877_ (.A1(_0544_),
    .A2(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3878_ (.A1(_0944_),
    .A2(_0949_),
    .B(_0952_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3879_ (.A1(_1811_),
    .A2(\Control_Unit.Q[1] ),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3880_ (.A1(_1800_),
    .A2(_1810_),
    .A3(\Control_Unit.Q[2] ),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3881_ (.A1(_0953_),
    .A2(_0954_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3882_ (.A1(_1799_),
    .A2(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3883_ (.A1(_1813_),
    .A2(_0544_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3884_ (.A1(_1926_),
    .A2(_0953_),
    .A3(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3885_ (.A1(_0958_),
    .A2(_0948_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3886_ (.A1(_0956_),
    .A2(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3887_ (.A1(_0956_),
    .A2(_0959_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3888_ (.A1(_0947_),
    .A2(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3889_ (.A1(_0542_),
    .A2(_0951_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3890_ (.A1(_0960_),
    .A2(_0962_),
    .B(_0963_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3891_ (.A1(_1810_),
    .A2(\Control_Unit.Q[2] ),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3892_ (.I(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3893_ (.A1(_1803_),
    .A2(\Control_Unit.Q[2] ),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3894_ (.A1(_1802_),
    .A2(_0965_),
    .A3(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3895_ (.A1(\Control_Unit.cont[1] ),
    .A2(_1770_),
    .A3(\Control_Unit.Q[3] ),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3896_ (.A1(_1796_),
    .A2(_0964_),
    .A3(_0968_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3897_ (.A1(_1820_),
    .A2(_0967_),
    .A3(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3898_ (.I(_1798_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3899_ (.A1(_0953_),
    .A2(_0954_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3900_ (.A1(_0971_),
    .A2(_0955_),
    .B(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3901_ (.A1(_0970_),
    .A2(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3902_ (.A1(_0961_),
    .A2(_0974_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3903_ (.I(_0946_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3904_ (.A1(_0961_),
    .A2(_0974_),
    .B(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3905_ (.A1(_0563_),
    .A2(_0951_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3906_ (.A1(_0975_),
    .A2(_0977_),
    .B(_0978_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3907_ (.I(_1910_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3908_ (.A1(_0965_),
    .A2(_0968_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3909_ (.A1(_0965_),
    .A2(_0968_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3910_ (.A1(_0971_),
    .A2(_0980_),
    .B(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3911_ (.A1(_1803_),
    .A2(_0557_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3912_ (.A1(_1811_),
    .A2(_0557_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3913_ (.A1(_0282_),
    .A2(_0983_),
    .B(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3914_ (.A1(_1800_),
    .A2(\Control_Unit.Q[4] ),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3915_ (.A1(_1933_),
    .A2(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3916_ (.A1(_1915_),
    .A2(_0985_),
    .A3(_0987_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3917_ (.A1(_0979_),
    .A2(_0982_),
    .A3(_0988_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3918_ (.A1(_1926_),
    .A2(_0965_),
    .A3(_0966_),
    .A4(_0969_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3919_ (.A1(_0967_),
    .A2(_0969_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3920_ (.A1(_1822_),
    .A2(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3921_ (.A1(_0990_),
    .A2(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3922_ (.A1(_0970_),
    .A2(_0973_),
    .B1(_0974_),
    .B2(_0961_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3923_ (.A1(_0989_),
    .A2(_0993_),
    .A3(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3924_ (.A1(_0586_),
    .A2(_0937_),
    .B1(_0940_),
    .B2(_0995_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3925_ (.I(_0939_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3926_ (.A1(_0982_),
    .A2(_0988_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3927_ (.A1(_0982_),
    .A2(_0988_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3928_ (.A1(_0979_),
    .A2(_0997_),
    .B(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3929_ (.A1(_0985_),
    .A2(_0987_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3930_ (.A1(_0985_),
    .A2(_0987_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3931_ (.A1(_1821_),
    .A2(_1000_),
    .B(_1001_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3932_ (.A1(_1801_),
    .A2(\Control_Unit.Q[4] ),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3933_ (.A1(_1797_),
    .A2(_0986_),
    .B(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3934_ (.A1(_1795_),
    .A2(\Control_Unit.Q[5] ),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3935_ (.A1(_1914_),
    .A2(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3936_ (.A1(_1004_),
    .A2(_1006_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3937_ (.A1(_0979_),
    .A2(_1007_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3938_ (.A1(_2070_),
    .A2(_1002_),
    .A3(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3939_ (.A1(_0990_),
    .A2(_0992_),
    .A3(_0989_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3940_ (.A1(_0990_),
    .A2(_0992_),
    .B(_0989_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3941_ (.A1(_1010_),
    .A2(_0994_),
    .B(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3942_ (.A1(_0999_),
    .A2(_1009_),
    .A3(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3943_ (.I(_0950_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3944_ (.A1(_0584_),
    .A2(_1014_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3945_ (.A1(_0996_),
    .A2(_1013_),
    .B(_1015_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3946_ (.A1(_0599_),
    .A2(_0951_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3947_ (.A1(_1004_),
    .A2(_1006_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3948_ (.A1(_2255_),
    .A2(_1007_),
    .B(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3949_ (.A1(_1796_),
    .A2(_0584_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3950_ (.A1(_1819_),
    .A2(_1005_),
    .B(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3951_ (.A1(_1769_),
    .A2(\Control_Unit.Q[6] ),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3952_ (.A1(_1785_),
    .A2(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3953_ (.A1(_1783_),
    .A2(_1020_),
    .A3(_1022_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3954_ (.A1(_1018_),
    .A2(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3955_ (.A1(_2067_),
    .A2(_1024_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3956_ (.A1(_1002_),
    .A2(_1008_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3957_ (.A1(_1002_),
    .A2(_1008_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3958_ (.A1(_0245_),
    .A2(_1026_),
    .B(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3959_ (.A1(_1025_),
    .A2(_1028_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3960_ (.A1(_0999_),
    .A2(_1009_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3961_ (.A1(_0999_),
    .A2(_1009_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3962_ (.A1(_1030_),
    .A2(_1012_),
    .B(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3963_ (.I(_0938_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3964_ (.A1(_1029_),
    .A2(_1032_),
    .B(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3965_ (.A1(_1029_),
    .A2(_1032_),
    .B(_1034_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3966_ (.A1(_1016_),
    .A2(_1035_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3967_ (.A1(_1018_),
    .A2(_1023_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3968_ (.A1(_0239_),
    .A2(_1024_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3969_ (.A1(_1020_),
    .A2(_1022_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3970_ (.A1(_1020_),
    .A2(_1022_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3971_ (.A1(_2070_),
    .A2(_1038_),
    .B(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3972_ (.A1(_1819_),
    .A2(_0599_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3973_ (.A1(_1825_),
    .A2(_1021_),
    .B(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3974_ (.A1(_1773_),
    .A2(\Control_Unit.Q[7] ),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3975_ (.A1(_1783_),
    .A2(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3976_ (.A1(_1848_),
    .A2(_1042_),
    .A3(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3977_ (.A1(_1040_),
    .A2(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3978_ (.A1(_0238_),
    .A2(_1046_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3979_ (.A1(_1036_),
    .A2(_1037_),
    .B(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3980_ (.A1(_1036_),
    .A2(_1037_),
    .A3(_1047_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3981_ (.A1(_1048_),
    .A2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3982_ (.A1(_1025_),
    .A2(_1028_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3983_ (.A1(_1029_),
    .A2(_1032_),
    .B(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3984_ (.A1(_1050_),
    .A2(_1052_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3985_ (.A1(_0611_),
    .A2(_1014_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3986_ (.A1(_0996_),
    .A2(_1053_),
    .B(_1054_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3987_ (.I(\Control_Unit.Q[8] ),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3988_ (.I(_1033_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3989_ (.A1(_1042_),
    .A2(_1044_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3990_ (.A1(_1042_),
    .A2(_1044_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3991_ (.A1(_1839_),
    .A2(_1057_),
    .B(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3992_ (.A1(_1824_),
    .A2(_0611_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3993_ (.A1(_1831_),
    .A2(_1043_),
    .B(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3994_ (.A1(\Control_Unit.cont[5] ),
    .A2(\Control_Unit.Q[8] ),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3995_ (.A1(_1776_),
    .A2(_1062_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3996_ (.A1(_1061_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3997_ (.A1(_0238_),
    .A2(_1064_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3998_ (.A1(_1059_),
    .A2(_1065_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3999_ (.A1(_2060_),
    .A2(_1066_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4000_ (.A1(_1040_),
    .A2(_1045_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4001_ (.A1(_1768_),
    .A2(_1046_),
    .B(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4002_ (.A1(_1067_),
    .A2(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4003_ (.A1(_1029_),
    .A2(_1032_),
    .B(_1048_),
    .C(_1051_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4004_ (.A1(_1049_),
    .A2(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4005_ (.A1(_1070_),
    .A2(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4006_ (.A1(_1055_),
    .A2(_0937_),
    .B1(_1056_),
    .B2(_1073_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4007_ (.I(\Control_Unit.Q[9] ),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4008_ (.A1(_1059_),
    .A2(_1065_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4009_ (.A1(_2112_),
    .A2(_1066_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4010_ (.I(_1061_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4011_ (.A1(_1766_),
    .A2(_1064_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4012_ (.A1(_1077_),
    .A2(_1063_),
    .B(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4013_ (.A1(_1838_),
    .A2(_1062_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4014_ (.A1(_1784_),
    .A2(_1055_),
    .B(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4015_ (.A1(_1776_),
    .A2(\Control_Unit.Q[9] ),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4016_ (.A1(_1765_),
    .A2(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4017_ (.A1(_1081_),
    .A2(_1083_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4018_ (.A1(_2059_),
    .A2(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4019_ (.A1(_0224_),
    .A2(_1079_),
    .A3(_1085_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4020_ (.A1(_1075_),
    .A2(_1076_),
    .B(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4021_ (.A1(_1075_),
    .A2(_1076_),
    .A3(_1086_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4022_ (.I(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4023_ (.A1(_1087_),
    .A2(_1089_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4024_ (.A1(_1067_),
    .A2(_1069_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4025_ (.A1(_1067_),
    .A2(_1069_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4026_ (.A1(_1091_),
    .A2(_1072_),
    .B(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4027_ (.A1(_1090_),
    .A2(_1093_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4028_ (.A1(_1074_),
    .A2(_0937_),
    .B1(_1056_),
    .B2(_1094_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4029_ (.A1(_1092_),
    .A2(_1087_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4030_ (.A1(_1049_),
    .A2(_1070_),
    .A3(_1071_),
    .B(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4031_ (.A1(_1081_),
    .A2(_1083_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4032_ (.A1(_2111_),
    .A2(_1084_),
    .B(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4033_ (.A1(_1765_),
    .A2(_1082_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4034_ (.A1(_1848_),
    .A2(_1074_),
    .B(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4035_ (.A1(_1760_),
    .A2(\Control_Unit.Q[10] ),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4036_ (.A1(_1752_),
    .A2(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4037_ (.A1(_1746_),
    .A2(_1100_),
    .A3(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4038_ (.A1(_0215_),
    .A2(_1098_),
    .A3(_1103_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4039_ (.A1(_1079_),
    .A2(_1085_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4040_ (.A1(_1079_),
    .A2(_1085_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4041_ (.A1(_2055_),
    .A2(_1105_),
    .B(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4042_ (.A1(_1104_),
    .A2(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4043_ (.A1(_1088_),
    .A2(_1096_),
    .B(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4044_ (.A1(_1088_),
    .A2(_1108_),
    .A3(_1096_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4045_ (.I(\Control_Unit.Mq ),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4046_ (.I(_1111_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4047_ (.I(\Control_Unit.Q[10] ),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4048_ (.A1(_1056_),
    .A2(_1109_),
    .A3(_1110_),
    .B1(_1112_),
    .B2(_1113_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4049_ (.I(\Control_Unit.Q[11] ),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4050_ (.I(_1111_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4051_ (.A1(_1104_),
    .A2(_1107_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4052_ (.A1(_1088_),
    .A2(_1108_),
    .A3(_1096_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4053_ (.A1(_1100_),
    .A2(_1102_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4054_ (.A1(_1100_),
    .A2(_1102_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4055_ (.A1(_1852_),
    .A2(_1118_),
    .B(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4056_ (.A1(_1752_),
    .A2(_1101_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4057_ (.A1(_1718_),
    .A2(_1113_),
    .B(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4058_ (.I(_1715_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4059_ (.A1(_1714_),
    .A2(\Control_Unit.Q[11] ),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4060_ (.A1(_1123_),
    .A2(_1124_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4061_ (.A1(_1857_),
    .A2(_1122_),
    .A3(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4062_ (.A1(_1120_),
    .A2(_1126_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4063_ (.A1(_0322_),
    .A2(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4064_ (.A1(_1098_),
    .A2(_1103_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4065_ (.A1(_1098_),
    .A2(_1103_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4066_ (.A1(_0222_),
    .A2(_1129_),
    .B(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4067_ (.A1(_1128_),
    .A2(_1131_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4068_ (.I(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4069_ (.A1(_1116_),
    .A2(_1117_),
    .B(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4070_ (.I(_1116_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4071_ (.I(_0946_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4072_ (.A1(_1135_),
    .A2(_1110_),
    .A3(_1132_),
    .B(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4073_ (.A1(_1114_),
    .A2(_1115_),
    .B1(_1134_),
    .B2(_1137_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4074_ (.A1(_1128_),
    .A2(_1131_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4075_ (.I(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4076_ (.A1(_1122_),
    .A2(_1125_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4077_ (.A1(_1122_),
    .A2(_1125_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4078_ (.A1(_2208_),
    .A2(_1140_),
    .B(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4079_ (.A1(_1123_),
    .A2(_1124_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4080_ (.A1(_2059_),
    .A2(_1114_),
    .B(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4081_ (.A1(_1715_),
    .A2(\Control_Unit.Q[12] ),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4082_ (.A1(_2046_),
    .A2(_1145_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4083_ (.A1(_0322_),
    .A2(_1144_),
    .A3(_1146_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4084_ (.A1(_1142_),
    .A2(_1147_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4085_ (.A1(_0351_),
    .A2(_1148_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4086_ (.A1(_1120_),
    .A2(_1126_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4087_ (.A1(_0317_),
    .A2(_1127_),
    .B(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4088_ (.A1(_1149_),
    .A2(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4089_ (.A1(_1139_),
    .A2(_1134_),
    .A3(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4090_ (.A1(_1135_),
    .A2(_1110_),
    .B(_1132_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4091_ (.I(_1152_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4092_ (.A1(_1138_),
    .A2(_1154_),
    .B(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4093_ (.I(\Control_Unit.Q[12] ),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4094_ (.A1(_0939_),
    .A2(_1153_),
    .A3(_1156_),
    .B1(_1112_),
    .B2(_1157_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4095_ (.I(\Control_Unit.Q[13] ),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4096_ (.A1(_1142_),
    .A2(_1147_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4097_ (.A1(_0320_),
    .A2(_1148_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4098_ (.A1(_1144_),
    .A2(_1146_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4099_ (.A1(_1144_),
    .A2(_1146_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4100_ (.A1(_2037_),
    .A2(_1161_),
    .B(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4101_ (.A1(_2047_),
    .A2(_1145_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4102_ (.A1(_0224_),
    .A2(_1157_),
    .B(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4103_ (.A1(_1716_),
    .A2(\Control_Unit.Q[13] ),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4104_ (.A1(_1868_),
    .A2(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4105_ (.A1(_0351_),
    .A2(_1165_),
    .A3(_1167_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4106_ (.A1(_1163_),
    .A2(_1168_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4107_ (.A1(_1889_),
    .A2(_1169_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4108_ (.A1(_1159_),
    .A2(_1160_),
    .B(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4109_ (.A1(_1159_),
    .A2(_1160_),
    .A3(_1170_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4110_ (.A1(_1171_),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4111_ (.A1(_1149_),
    .A2(_1151_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4112_ (.A1(_1174_),
    .A2(_1156_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4113_ (.A1(_1173_),
    .A2(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4114_ (.A1(_1158_),
    .A2(_1115_),
    .B1(_1056_),
    .B2(_1176_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4115_ (.I(\Control_Unit.Q[14] ),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4116_ (.A1(_1139_),
    .A2(_1134_),
    .B(_1152_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4117_ (.A1(_1174_),
    .A2(_1171_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4118_ (.A1(_1165_),
    .A2(_1167_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4119_ (.A1(_1165_),
    .A2(_1167_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4120_ (.A1(_0319_),
    .A2(_1180_),
    .B(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4121_ (.A1(_1868_),
    .A2(_1166_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4122_ (.A1(_0215_),
    .A2(_1158_),
    .B(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4123_ (.A1(\Control_Unit.cont[11] ),
    .A2(\Control_Unit.Q[14] ),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4124_ (.A1(_1711_),
    .A2(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4125_ (.A1(_1735_),
    .A2(_1184_),
    .A3(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4126_ (.A1(_1182_),
    .A2(_1187_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4127_ (.A1(_0388_),
    .A2(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4128_ (.A1(_1163_),
    .A2(_1168_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4129_ (.A1(_1882_),
    .A2(_1169_),
    .B(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4130_ (.A1(_1189_),
    .A2(_1191_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4131_ (.I(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4132_ (.A1(_1178_),
    .A2(_1179_),
    .B(_1193_),
    .C(_1172_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4133_ (.A1(_1178_),
    .A2(_1179_),
    .B(_1172_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4134_ (.A1(_1192_),
    .A2(_1195_),
    .B(_0976_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4135_ (.A1(_1177_),
    .A2(_1115_),
    .B1(_1194_),
    .B2(_1196_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4136_ (.A1(_1182_),
    .A2(_1187_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4137_ (.A1(_2177_),
    .A2(_1188_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4138_ (.A1(_1184_),
    .A2(_1186_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4139_ (.A1(_1184_),
    .A2(_1186_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4140_ (.A1(_1879_),
    .A2(_1199_),
    .B(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4141_ (.A1(_1736_),
    .A2(_1185_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4142_ (.A1(_1713_),
    .A2(_1177_),
    .B(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4143_ (.A1(\Control_Unit.cont[12] ),
    .A2(\Control_Unit.Q[15] ),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4144_ (.A1(_1712_),
    .A2(_1204_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4145_ (.A1(_1203_),
    .A2(_1205_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4146_ (.A1(_1710_),
    .A2(_1206_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4147_ (.A1(_1201_),
    .A2(_1207_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4148_ (.A1(_0383_),
    .A2(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4149_ (.A1(_1197_),
    .A2(_1198_),
    .B(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4150_ (.A1(_1197_),
    .A2(_1198_),
    .A3(_1209_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4151_ (.A1(_1210_),
    .A2(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4152_ (.A1(_1189_),
    .A2(_1191_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4153_ (.A1(_1213_),
    .A2(_1194_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4154_ (.A1(_1212_),
    .A2(_1214_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4155_ (.A1(_0714_),
    .A2(_1014_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4156_ (.A1(_0996_),
    .A2(_1215_),
    .B(_1216_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4157_ (.A1(_1736_),
    .A2(_0714_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4158_ (.A1(_1712_),
    .A2(_1204_),
    .B(_1217_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4159_ (.A1(\Control_Unit.cont[13] ),
    .A2(\Control_Unit.Q[16] ),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4160_ (.A1(_1709_),
    .A2(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4161_ (.A1(_1218_),
    .A2(_1220_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4162_ (.A1(_1706_),
    .A2(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4163_ (.A1(_1203_),
    .A2(_1205_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4164_ (.A1(_2027_),
    .A2(_1206_),
    .B(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4165_ (.A1(_1222_),
    .A2(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4166_ (.A1(_1201_),
    .A2(_1207_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4167_ (.A1(_0383_),
    .A2(_1208_),
    .B(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4168_ (.A1(_1225_),
    .A2(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4169_ (.A1(_1213_),
    .A2(_1210_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4170_ (.I(_1211_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4171_ (.A1(_1194_),
    .A2(_1229_),
    .B(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4172_ (.A1(_1228_),
    .A2(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4173_ (.A1(_1228_),
    .A2(_1231_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4174_ (.I(\Control_Unit.Q[16] ),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4175_ (.A1(_0939_),
    .A2(_1232_),
    .A3(_1233_),
    .B1(_0936_),
    .B2(_1234_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4176_ (.A1(_1225_),
    .A2(_1227_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4177_ (.A1(_1235_),
    .A2(_1233_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4178_ (.A1(_1222_),
    .A2(_1224_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4179_ (.A1(_1734_),
    .A2(\Control_Unit.Q[17] ),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4180_ (.A1(\Control_Unit.cont[15] ),
    .A2(_1238_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4181_ (.A1(_1735_),
    .A2(_1234_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4182_ (.A1(_1734_),
    .A2(_1219_),
    .B(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4183_ (.A1(_1239_),
    .A2(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4184_ (.A1(_1218_),
    .A2(_1220_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4185_ (.A1(_1728_),
    .A2(_1221_),
    .B(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4186_ (.A1(_1242_),
    .A2(_1244_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4187_ (.A1(_1242_),
    .A2(_1244_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4188_ (.A1(_1245_),
    .A2(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4189_ (.A1(_1237_),
    .A2(_1247_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4190_ (.A1(_1236_),
    .A2(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4191_ (.A1(_0743_),
    .A2(_1014_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4192_ (.A1(_0996_),
    .A2(_1249_),
    .B(_1250_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4193_ (.I(\Control_Unit.Q[18] ),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4194_ (.A1(_1237_),
    .A2(_1235_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4195_ (.A1(_1228_),
    .A2(_1248_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4196_ (.A1(_1247_),
    .A2(_1252_),
    .B1(_1253_),
    .B2(_1231_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4197_ (.A1(_1706_),
    .A2(_1251_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4198_ (.A1(_2026_),
    .A2(_0743_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4199_ (.A1(_1706_),
    .A2(_1238_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4200_ (.A1(_1256_),
    .A2(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4201_ (.A1(_1255_),
    .A2(_1258_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4202_ (.I(_1241_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4203_ (.A1(_1239_),
    .A2(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4204_ (.A1(_1261_),
    .A2(_1245_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4205_ (.A1(_1259_),
    .A2(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4206_ (.A1(_1254_),
    .A2(_1263_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4207_ (.A1(_1254_),
    .A2(_1263_),
    .B(_1136_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4208_ (.A1(_1251_),
    .A2(_1115_),
    .B1(_1264_),
    .B2(_1265_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4209_ (.A1(_1261_),
    .A2(_1259_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4210_ (.A1(_1256_),
    .A2(_1257_),
    .B(_1255_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4211_ (.A1(_1707_),
    .A2(_0768_),
    .B(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4212_ (.A1(\Control_Unit.Q[19] ),
    .A2(_1268_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4213_ (.I(_1269_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4214_ (.A1(_1245_),
    .A2(_1259_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4215_ (.A1(_1264_),
    .A2(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4216_ (.A1(_1266_),
    .A2(_1270_),
    .A3(_1272_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4217_ (.I(_0950_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4218_ (.A1(_0788_),
    .A2(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4219_ (.A1(_0940_),
    .A2(_1273_),
    .B(_1275_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4220_ (.A1(_1263_),
    .A2(_1270_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4221_ (.A1(_1247_),
    .A2(_1252_),
    .A3(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4222_ (.A1(_1261_),
    .A2(_1269_),
    .B(_1259_),
    .C(_1245_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4223_ (.A1(_1266_),
    .A2(_1270_),
    .B(_1277_),
    .C(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4224_ (.A1(_1253_),
    .A2(_1276_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4225_ (.I(_1280_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4226_ (.A1(_1194_),
    .A2(_1229_),
    .B(_1281_),
    .C(_1230_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4227_ (.A1(_0788_),
    .A2(_1267_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4228_ (.A1(_0383_),
    .A2(_0768_),
    .A3(\Control_Unit.Q[19] ),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4229_ (.A1(_0797_),
    .A2(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4230_ (.A1(_1283_),
    .A2(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4231_ (.A1(_1279_),
    .A2(_1282_),
    .B(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4232_ (.A1(_1286_),
    .A2(_1279_),
    .A3(_1282_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4233_ (.A1(_0947_),
    .A2(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4234_ (.A1(_0797_),
    .A2(_1274_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4235_ (.A1(_1287_),
    .A2(_1289_),
    .B(_1290_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4236_ (.A1(_1283_),
    .A2(_1285_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4237_ (.A1(_1291_),
    .A2(_1287_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4238_ (.A1(_1708_),
    .A2(_0768_),
    .A3(_0788_),
    .A4(_0797_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4239_ (.A1(_0814_),
    .A2(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4240_ (.A1(_1292_),
    .A2(_1294_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4241_ (.A1(_0814_),
    .A2(_1274_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4242_ (.A1(_0940_),
    .A2(_1295_),
    .B(_1296_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4243_ (.I(_0822_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4244_ (.A1(_1283_),
    .A2(_1285_),
    .B(_1293_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4245_ (.A1(_0814_),
    .A2(_1298_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4246_ (.A1(_1287_),
    .A2(_1294_),
    .B(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4247_ (.A1(_1297_),
    .A2(_1300_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4248_ (.A1(_1297_),
    .A2(_1300_),
    .B(_1136_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4249_ (.A1(_1297_),
    .A2(_1112_),
    .B1(_1301_),
    .B2(_1302_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4250_ (.A1(_1297_),
    .A2(_1033_),
    .A3(_1300_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4251_ (.A1(_0936_),
    .A2(_1302_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4252_ (.I0(_1303_),
    .I1(_1304_),
    .S(_0841_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4253_ (.I(_1305_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4254_ (.I(\Control_Unit.Q[24] ),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4255_ (.A1(_1174_),
    .A2(_1171_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4256_ (.I(_1172_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4257_ (.A1(_1156_),
    .A2(_1307_),
    .B(_1192_),
    .C(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4258_ (.I(_1229_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4259_ (.A1(_1309_),
    .A2(_1310_),
    .B(_1280_),
    .C(_1211_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4260_ (.A1(_0822_),
    .A2(_0841_),
    .A3(_1294_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4261_ (.A1(_1286_),
    .A2(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4262_ (.A1(_0822_),
    .A2(_0841_),
    .A3(_1299_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4263_ (.A1(_1286_),
    .A2(_1279_),
    .A3(_1312_),
    .B(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4264_ (.A1(_1311_),
    .A2(_1313_),
    .B(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4265_ (.A1(_0938_),
    .A2(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4266_ (.I(_1306_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4267_ (.A1(_1318_),
    .A2(_1316_),
    .B(_1136_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4268_ (.A1(_1111_),
    .A2(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4269_ (.A1(_1306_),
    .A2(_1317_),
    .B(_1320_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4270_ (.I(_1321_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4271_ (.I(\Control_Unit.Q[25] ),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4272_ (.A1(_1306_),
    .A2(_1317_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4273_ (.A1(_1322_),
    .A2(_1320_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4274_ (.A1(_1322_),
    .A2(_1323_),
    .B(_1324_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4275_ (.A1(\Control_Unit.Q[24] ),
    .A2(_1322_),
    .A3(\Control_Unit.Q[26] ),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4276_ (.A1(_1316_),
    .A2(_1325_),
    .B(_0946_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4277_ (.A1(_1306_),
    .A2(_1322_),
    .A3(_1317_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4278_ (.I(\Control_Unit.Q[26] ),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4279_ (.A1(_1112_),
    .A2(_1326_),
    .B1(_1327_),
    .B2(_1328_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4280_ (.A1(_1111_),
    .A2(_1326_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4281_ (.A1(_0895_),
    .A2(_1325_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4282_ (.A1(_0895_),
    .A2(_1329_),
    .B1(_1330_),
    .B2(_1317_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4283_ (.I(_1331_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4284_ (.I(\Control_Unit.Q[28] ),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4285_ (.I(_0895_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4286_ (.A1(_1333_),
    .A2(_1316_),
    .A3(_1325_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4287_ (.I(_1334_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4288_ (.A1(_1332_),
    .A2(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4289_ (.A1(_0490_),
    .A2(_1336_),
    .B(_0950_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4290_ (.A1(_0947_),
    .A2(_1335_),
    .B(_1332_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4291_ (.A1(_1337_),
    .A2(_1338_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4292_ (.I(\Control_Unit.Q[29] ),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4293_ (.A1(_1332_),
    .A2(_1339_),
    .A3(_0976_),
    .A4(_1335_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4294_ (.A1(_1339_),
    .A2(_1337_),
    .B(_1340_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4295_ (.A1(_1332_),
    .A2(\Control_Unit.Q[29] ),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4296_ (.A1(_1335_),
    .A2(_1341_),
    .B(_0927_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4297_ (.A1(_0927_),
    .A2(_1334_),
    .A3(_1341_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4298_ (.A1(_1033_),
    .A2(_1343_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4299_ (.A1(_0927_),
    .A2(_1274_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4300_ (.A1(_1342_),
    .A2(_1344_),
    .B(_1345_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4301_ (.A1(\Control_Unit.Q[31] ),
    .A2(_0936_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4302_ (.A1(_0976_),
    .A2(_1343_),
    .B(\Control_Unit.Q[31] ),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4303_ (.A1(_1344_),
    .A2(_1346_),
    .B(_1347_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4304_ (.A1(_0338_),
    .A2(\Control_Unit.Mc ),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4305_ (.I(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4306_ (.I(_1349_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4307_ (.A1(_0525_),
    .A2(_0941_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4308_ (.I(\Control_Unit.Mc ),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4309_ (.I(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4310_ (.I(_1353_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4311_ (.A1(_0525_),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4312_ (.A1(_1350_),
    .A2(_1351_),
    .B(_1355_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4313_ (.I(_1348_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4314_ (.I(_1356_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4315_ (.A1(\Control_Unit.C[1] ),
    .A2(_0282_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4316_ (.I(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4317_ (.I(_2013_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4318_ (.A1(_1360_),
    .A2(_1809_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4319_ (.A1(_0525_),
    .A2(_0941_),
    .B1(_1359_),
    .B2(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4320_ (.A1(_2014_),
    .A2(_2153_),
    .A3(_1359_),
    .A4(_1361_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4321_ (.I(\Control_Unit.Mc ),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4322_ (.I(_1364_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4323_ (.A1(_1357_),
    .A2(_1362_),
    .A3(_1363_),
    .B1(_1365_),
    .B2(_1360_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4324_ (.A1(\Control_Unit.C[2] ),
    .A2(_1795_),
    .A3(_1803_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4325_ (.A1(_1358_),
    .A2(_1366_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4326_ (.A1(_1359_),
    .A2(_1366_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4327_ (.A1(_1367_),
    .A2(_1368_),
    .B(_1363_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4328_ (.A1(\Control_Unit.C[0] ),
    .A2(_1814_),
    .A3(_1359_),
    .A4(_1361_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4329_ (.A1(_1370_),
    .A2(_1366_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4330_ (.A1(_1357_),
    .A2(_1369_),
    .A3(_1371_),
    .B1(_1365_),
    .B2(_0541_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4331_ (.A1(_2015_),
    .A2(_1354_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4332_ (.A1(_1915_),
    .A2(\Control_Unit.C[3] ),
    .A3(_1802_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4333_ (.A1(\Control_Unit.C[2] ),
    .A2(_1804_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4334_ (.A1(_2016_),
    .A2(_1804_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4335_ (.A1(_1798_),
    .A2(_1374_),
    .B(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4336_ (.A1(_1373_),
    .A2(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4337_ (.A1(_1367_),
    .A2(_1377_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4338_ (.I(_1348_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4339_ (.A1(_1371_),
    .A2(_1378_),
    .B(_1379_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4340_ (.A1(_1371_),
    .A2(_1378_),
    .B(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4341_ (.A1(_1372_),
    .A2(_1381_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4342_ (.A1(_1373_),
    .A2(_1376_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4343_ (.A1(_1825_),
    .A2(\Control_Unit.C[4] ),
    .A3(_1797_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4344_ (.A1(\Control_Unit.C[3] ),
    .A2(_1807_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4345_ (.A1(_2015_),
    .A2(_1807_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4346_ (.A1(_1915_),
    .A2(_1384_),
    .B(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4347_ (.A1(_1383_),
    .A2(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4348_ (.A1(_1382_),
    .A2(_1387_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4349_ (.A1(_1367_),
    .A2(_1373_),
    .A3(_1376_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4350_ (.A1(_1370_),
    .A2(_1366_),
    .A3(_1389_),
    .B1(_1377_),
    .B2(_1367_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4351_ (.A1(_1388_),
    .A2(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4352_ (.A1(_2009_),
    .A2(_1354_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4353_ (.A1(_1350_),
    .A2(_1391_),
    .B(_1392_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4354_ (.A1(_1383_),
    .A2(_1386_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4355_ (.I(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4356_ (.A1(_1382_),
    .A2(_1387_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4357_ (.A1(_1388_),
    .A2(_1390_),
    .B(_1395_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4358_ (.A1(_1831_),
    .A2(_1820_),
    .A3(_2006_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4359_ (.A1(_2008_),
    .A2(_0971_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4360_ (.A1(_2008_),
    .A2(_0971_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4361_ (.A1(_0979_),
    .A2(_1398_),
    .B(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4362_ (.A1(_1397_),
    .A2(_1400_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4363_ (.A1(_1394_),
    .A2(_1396_),
    .A3(_1401_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4364_ (.I(_1352_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4365_ (.A1(_2007_),
    .A2(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4366_ (.A1(_1350_),
    .A2(_1402_),
    .B(_1404_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4367_ (.I(_2011_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4368_ (.I(\Control_Unit.Mc ),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4369_ (.I(_1406_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4370_ (.A1(_1394_),
    .A2(_1401_),
    .B(_1390_),
    .C(_1388_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4371_ (.A1(_1394_),
    .A2(_1395_),
    .B(_1401_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4372_ (.A1(_1408_),
    .A2(_1409_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4373_ (.A1(_1397_),
    .A2(_1400_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4374_ (.A1(_1824_),
    .A2(\Control_Unit.C[6] ),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4375_ (.A1(_1838_),
    .A2(_1412_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4376_ (.A1(_2073_),
    .A2(\Control_Unit.C[5] ),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4377_ (.A1(_2073_),
    .A2(_2006_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4378_ (.A1(_1784_),
    .A2(_1414_),
    .B(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4379_ (.A1(_1413_),
    .A2(_1416_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4380_ (.A1(_1411_),
    .A2(_1417_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4381_ (.A1(_1410_),
    .A2(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4382_ (.A1(_0421_),
    .A2(_1352_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4383_ (.I(_1420_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4384_ (.I(_1421_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4385_ (.A1(_1410_),
    .A2(_1418_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4386_ (.A1(_1422_),
    .A2(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4387_ (.A1(_1405_),
    .A2(_1407_),
    .B1(_1419_),
    .B2(_1424_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4388_ (.A1(_1411_),
    .A2(_1417_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4389_ (.A1(_1425_),
    .A2(_1423_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4390_ (.A1(_1413_),
    .A2(_1416_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4391_ (.A1(_1839_),
    .A2(_1412_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4392_ (.A1(_1910_),
    .A2(_1405_),
    .B(_1428_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4393_ (.A1(_1831_),
    .A2(\Control_Unit.C[7] ),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4394_ (.A1(_1765_),
    .A2(_1430_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4395_ (.A1(_1429_),
    .A2(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4396_ (.A1(_1427_),
    .A2(_1432_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4397_ (.A1(_1426_),
    .A2(_1433_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4398_ (.A1(_2010_),
    .A2(_1403_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4399_ (.A1(_1350_),
    .A2(_1434_),
    .B(_1435_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4400_ (.I(_1356_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4401_ (.I(_1418_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4402_ (.A1(_1408_),
    .A2(_1409_),
    .B(_1437_),
    .C(_1433_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4403_ (.I(_1432_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4404_ (.A1(_1427_),
    .A2(_1425_),
    .B(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4405_ (.A1(_1438_),
    .A2(_1440_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4406_ (.A1(_1429_),
    .A2(_1431_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4407_ (.A1(_1838_),
    .A2(\Control_Unit.C[8] ),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4408_ (.A1(_2059_),
    .A2(_1443_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4409_ (.A1(_1832_),
    .A2(\Control_Unit.C[7] ),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4410_ (.A1(_1766_),
    .A2(_1430_),
    .B(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4411_ (.A1(_1444_),
    .A2(_1446_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4412_ (.A1(_1444_),
    .A2(_1446_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4413_ (.A1(_1447_),
    .A2(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4414_ (.A1(_1442_),
    .A2(_1449_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4415_ (.A1(_1441_),
    .A2(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4416_ (.A1(_2001_),
    .A2(_1407_),
    .B1(_1436_),
    .B2(_1451_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4417_ (.A1(_1442_),
    .A2(_1449_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4418_ (.I(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4419_ (.A1(_1441_),
    .A2(_1450_),
    .B(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4420_ (.A1(_1760_),
    .A2(\Control_Unit.C[9] ),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4421_ (.A1(_1123_),
    .A2(_1455_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4422_ (.A1(_1759_),
    .A2(_1443_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4423_ (.A1(_2067_),
    .A2(_2001_),
    .B(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4424_ (.A1(_1456_),
    .A2(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4425_ (.A1(_1447_),
    .A2(_1459_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4426_ (.A1(_1454_),
    .A2(_1460_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4427_ (.A1(_2000_),
    .A2(_1407_),
    .B1(_1436_),
    .B2(_1461_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4428_ (.I(_1364_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4429_ (.A1(_1438_),
    .A2(_1440_),
    .B(_1450_),
    .C(_1460_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4430_ (.A1(_1447_),
    .A2(_1452_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4431_ (.A1(_1459_),
    .A2(_1464_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4432_ (.A1(_1456_),
    .A2(_1458_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4433_ (.A1(_1752_),
    .A2(\Control_Unit.C[10] ),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4434_ (.A1(_2046_),
    .A2(_1467_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4435_ (.A1(_1852_),
    .A2(_1455_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4436_ (.A1(_0238_),
    .A2(_2000_),
    .B(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4437_ (.A1(_1468_),
    .A2(_1470_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4438_ (.A1(_1466_),
    .A2(_1471_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4439_ (.I(_1472_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4440_ (.A1(_1463_),
    .A2(_1465_),
    .B(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4441_ (.A1(_1463_),
    .A2(_1465_),
    .A3(_1473_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4442_ (.A1(_1422_),
    .A2(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4443_ (.A1(_2004_),
    .A2(_1462_),
    .B1(_1474_),
    .B2(_1476_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4444_ (.A1(_1466_),
    .A2(_1471_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4445_ (.I(_1477_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4446_ (.A1(_1478_),
    .A2(_1474_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4447_ (.A1(_1468_),
    .A2(_1470_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4448_ (.A1(_1123_),
    .A2(\Control_Unit.C[11] ),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4449_ (.A1(_2036_),
    .A2(_1481_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4450_ (.A1(_2047_),
    .A2(_1467_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4451_ (.A1(_2060_),
    .A2(_2004_),
    .B(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4452_ (.A1(_1482_),
    .A2(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4453_ (.A1(_1480_),
    .A2(_1485_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4454_ (.A1(_1479_),
    .A2(_1486_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4455_ (.A1(_1479_),
    .A2(_1486_),
    .B(_1421_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4456_ (.A1(_2003_),
    .A2(_1462_),
    .B1(_1487_),
    .B2(_1488_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4457_ (.A1(_1480_),
    .A2(_1485_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4458_ (.A1(_1482_),
    .A2(_1484_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4459_ (.A1(_2046_),
    .A2(\Control_Unit.C[12] ),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4460_ (.A1(_2041_),
    .A2(_1491_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4461_ (.A1(_2036_),
    .A2(_1481_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4462_ (.A1(_0224_),
    .A2(_2003_),
    .B(_1493_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4463_ (.A1(_1492_),
    .A2(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4464_ (.A1(_1490_),
    .A2(_1495_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4465_ (.A1(_1489_),
    .A2(_1487_),
    .A3(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4466_ (.I(_1489_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4467_ (.A1(_1478_),
    .A2(_1474_),
    .B(_1486_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4468_ (.I(_1496_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4469_ (.A1(_1498_),
    .A2(_1499_),
    .B(_1500_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4470_ (.I(_2019_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4471_ (.A1(_1349_),
    .A2(_1497_),
    .A3(_1501_),
    .B1(_1365_),
    .B2(_1502_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4472_ (.I(_2018_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4473_ (.A1(_1490_),
    .A2(_1495_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4474_ (.I(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4475_ (.A1(_1492_),
    .A2(_1494_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4476_ (.A1(_2036_),
    .A2(\Control_Unit.C[13] ),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4477_ (.A1(_1879_),
    .A2(_1507_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4478_ (.A1(_0319_),
    .A2(_1491_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4479_ (.A1(_0215_),
    .A2(_1502_),
    .B(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4480_ (.A1(_1508_),
    .A2(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4481_ (.A1(_1506_),
    .A2(_1511_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4482_ (.A1(_1505_),
    .A2(_1501_),
    .A3(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4483_ (.I(_1420_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4484_ (.A1(_1505_),
    .A2(_1501_),
    .B(_1512_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4485_ (.A1(_1514_),
    .A2(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4486_ (.A1(_1503_),
    .A2(_1462_),
    .B1(_1513_),
    .B2(_1516_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4487_ (.A1(_1506_),
    .A2(_1511_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4488_ (.A1(_1508_),
    .A2(_1510_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4489_ (.A1(_2041_),
    .A2(\Control_Unit.C[14] ),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4490_ (.A1(_2026_),
    .A2(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4491_ (.A1(_1880_),
    .A2(_1507_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4492_ (.A1(_0322_),
    .A2(_1503_),
    .B(_1521_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4493_ (.A1(_1520_),
    .A2(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4494_ (.A1(_1518_),
    .A2(_1523_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4495_ (.I(_1524_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4496_ (.A1(_1517_),
    .A2(_1515_),
    .A3(_1525_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4497_ (.A1(_1517_),
    .A2(_1515_),
    .B(_1525_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4498_ (.I(_2021_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4499_ (.A1(_1349_),
    .A2(_1526_),
    .A3(_1527_),
    .B1(_1406_),
    .B2(_1528_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4500_ (.A1(_1518_),
    .A2(_1523_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4501_ (.I(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4502_ (.A1(_1520_),
    .A2(_1522_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4503_ (.A1(_2027_),
    .A2(_1519_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4504_ (.A1(_0351_),
    .A2(_1528_),
    .B(_1532_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4505_ (.A1(_1879_),
    .A2(\Control_Unit.C[15] ),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4506_ (.A1(_1707_),
    .A2(_1534_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4507_ (.A1(_1533_),
    .A2(_1535_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4508_ (.A1(_1531_),
    .A2(_1536_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4509_ (.A1(_1530_),
    .A2(_1527_),
    .A3(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4510_ (.A1(_1530_),
    .A2(_1527_),
    .B(_1537_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4511_ (.A1(_1422_),
    .A2(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4512_ (.A1(_2020_),
    .A2(_1403_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4513_ (.A1(_1538_),
    .A2(_1540_),
    .B(_1541_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4514_ (.I(_1989_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4515_ (.A1(_1531_),
    .A2(_1536_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4516_ (.A1(_1543_),
    .A2(_1539_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4517_ (.A1(_2026_),
    .A2(\Control_Unit.C[16] ),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4518_ (.A1(_1880_),
    .A2(\Control_Unit.C[15] ),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4519_ (.A1(_1728_),
    .A2(_1534_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4520_ (.A1(_1546_),
    .A2(_1547_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4521_ (.A1(_1545_),
    .A2(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4522_ (.A1(_1533_),
    .A2(_1535_),
    .A3(_1549_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4523_ (.I(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4524_ (.A1(_1533_),
    .A2(_1535_),
    .B(_1549_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4525_ (.A1(_1551_),
    .A2(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4526_ (.A1(_1544_),
    .A2(_1553_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4527_ (.A1(_1544_),
    .A2(_1553_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4528_ (.A1(_1514_),
    .A2(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4529_ (.A1(_1542_),
    .A2(_1462_),
    .B1(_1554_),
    .B2(_1556_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4530_ (.A1(_1988_),
    .A2(_1354_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4531_ (.A1(_1550_),
    .A2(_1555_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4532_ (.A1(_1728_),
    .A2(_1987_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4533_ (.A1(_1546_),
    .A2(_1547_),
    .B(_1545_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4534_ (.A1(_0388_),
    .A2(_1542_),
    .B(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4535_ (.A1(_1559_),
    .A2(_1561_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4536_ (.A1(_1558_),
    .A2(_1562_),
    .B(_1379_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4537_ (.A1(_1558_),
    .A2(_1562_),
    .B(_1563_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4538_ (.A1(_1557_),
    .A2(_1564_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4539_ (.I(_1992_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4540_ (.A1(_1544_),
    .A2(_1553_),
    .B(_1551_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4541_ (.I(_1562_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4542_ (.A1(_1546_),
    .A2(_1547_),
    .B(_1545_),
    .C(_1559_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4543_ (.A1(_1566_),
    .A2(_1567_),
    .B(_1568_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4544_ (.A1(_2176_),
    .A2(_1989_),
    .A3(_1559_),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4545_ (.A1(_1708_),
    .A2(_1988_),
    .B(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4546_ (.A1(_1565_),
    .A2(_1571_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4547_ (.A1(_1569_),
    .A2(_1572_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4548_ (.A1(_1569_),
    .A2(_1572_),
    .B(_1421_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4549_ (.A1(_1565_),
    .A2(_1365_),
    .B1(_1573_),
    .B2(_1574_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4550_ (.A1(_1993_),
    .A2(_1570_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4551_ (.A1(_1569_),
    .A2(_1572_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4552_ (.A1(_0384_),
    .A2(_1988_),
    .A3(_1993_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4553_ (.A1(_1991_),
    .A2(_1577_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4554_ (.A1(_1990_),
    .A2(_1577_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4555_ (.A1(_1575_),
    .A2(_1576_),
    .B(_1578_),
    .C(_1579_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4556_ (.A1(_1578_),
    .A2(_1579_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4557_ (.A1(_1993_),
    .A2(_1570_),
    .B(_1573_),
    .C(_1581_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4558_ (.I(_1991_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4559_ (.A1(_1349_),
    .A2(_1580_),
    .A3(_1582_),
    .B1(_1406_),
    .B2(_1583_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4560_ (.I(_1983_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4561_ (.A1(_1991_),
    .A2(_1572_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4562_ (.A1(_1550_),
    .A2(_1567_),
    .B(_1568_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4563_ (.A1(_1585_),
    .A2(_1586_),
    .B(_1579_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4564_ (.A1(_1575_),
    .A2(_1578_),
    .B(_1587_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4565_ (.A1(_1553_),
    .A2(_1562_),
    .A3(_1585_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4566_ (.A1(_1543_),
    .A2(_1539_),
    .B(_1589_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4567_ (.A1(_1588_),
    .A2(_1590_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4568_ (.A1(_1588_),
    .A2(_1590_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4569_ (.A1(_1584_),
    .A2(_1592_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4570_ (.A1(_0421_),
    .A2(_1593_),
    .B(_1364_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4571_ (.A1(_1584_),
    .A2(_1594_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4572_ (.A1(_1584_),
    .A2(_1436_),
    .A3(_1591_),
    .B(_1595_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4573_ (.A1(_1422_),
    .A2(_1593_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4574_ (.A1(_1982_),
    .A2(_1594_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4575_ (.A1(_1982_),
    .A2(_1596_),
    .B(_1597_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4576_ (.A1(_1982_),
    .A2(_1593_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4577_ (.A1(_1981_),
    .A2(_1985_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4578_ (.A1(_1584_),
    .A2(_1592_),
    .A3(_1599_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4579_ (.A1(_0421_),
    .A2(_1600_),
    .B(_1364_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4580_ (.A1(_1985_),
    .A2(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4581_ (.A1(_1985_),
    .A2(_1436_),
    .A3(_1598_),
    .B(_1602_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4582_ (.I(_1984_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4583_ (.A1(_1588_),
    .A2(_1590_),
    .B(_1599_),
    .C(_1983_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(_1603_),
    .A2(_1601_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4585_ (.A1(_1603_),
    .A2(_1357_),
    .A3(_1604_),
    .B(_1605_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4586_ (.I(_1977_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4587_ (.I(_1603_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4588_ (.A1(_1607_),
    .A2(_1606_),
    .A3(_1604_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4589_ (.A1(_1356_),
    .A2(_1608_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4590_ (.A1(_1353_),
    .A2(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4591_ (.A1(_1603_),
    .A2(_1600_),
    .A3(_1609_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4592_ (.A1(_1606_),
    .A2(_1610_),
    .B(_1611_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4593_ (.I(_1976_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4594_ (.A1(_1421_),
    .A2(_1608_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4595_ (.A1(_1612_),
    .A2(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4596_ (.A1(_1612_),
    .A2(_1610_),
    .B(_1614_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4597_ (.A1(_1612_),
    .A2(_1979_),
    .A3(_1608_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4598_ (.A1(_0490_),
    .A2(_1615_),
    .B(_1353_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4599_ (.A1(_1612_),
    .A2(_1613_),
    .B(_1979_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4600_ (.A1(_1616_),
    .A2(_1617_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4601_ (.I(_1978_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4602_ (.A1(_1978_),
    .A2(_1379_),
    .A3(_1615_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4603_ (.A1(_1618_),
    .A2(_1616_),
    .B(_1619_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4604_ (.I(_1996_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4605_ (.A1(_1976_),
    .A2(_1978_),
    .A3(_1979_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4606_ (.A1(_1607_),
    .A2(_1606_),
    .A3(_1604_),
    .A4(_1621_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4607_ (.I(_1622_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4608_ (.A1(_1620_),
    .A2(_1623_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4609_ (.A1(_0490_),
    .A2(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4610_ (.A1(_1514_),
    .A2(_1623_),
    .B(_1620_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4611_ (.A1(_1407_),
    .A2(_1625_),
    .B(_1626_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4612_ (.I(_1995_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4613_ (.A1(_1620_),
    .A2(_1623_),
    .B(_1356_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4614_ (.A1(_1353_),
    .A2(_1628_),
    .B(_1627_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4615_ (.A1(_1627_),
    .A2(_1357_),
    .A3(_1624_),
    .B(_1629_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4616_ (.I(_1997_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4617_ (.A1(_1627_),
    .A2(_1620_),
    .A3(_1623_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(_1997_),
    .A2(_1403_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4619_ (.A1(_1627_),
    .A2(_1996_),
    .A3(_1997_),
    .A4(_1622_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4620_ (.A1(_1379_),
    .A2(_1633_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4621_ (.A1(_1630_),
    .A2(_1631_),
    .B1(_1632_),
    .B2(_1634_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4622_ (.A1(\Control_Unit.C[31] ),
    .A2(_1406_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4623_ (.A1(_1514_),
    .A2(_1633_),
    .B(\Control_Unit.C[31] ),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4624_ (.A1(_1634_),
    .A2(_1635_),
    .B(_1636_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4625_ (.A1(_0941_),
    .A2(_0532_),
    .B(_0340_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4626_ (.A1(_0506_),
    .A2(_0532_),
    .B(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4627_ (.A1(_0533_),
    .A2(_0363_),
    .B(_1638_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4628_ (.A1(_0506_),
    .A2(_0532_),
    .B(_0280_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4629_ (.I(_0377_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4630_ (.A1(_0281_),
    .A2(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4631_ (.I(_0375_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4632_ (.A1(_0536_),
    .A2(_1642_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4633_ (.A1(_1639_),
    .A2(_1641_),
    .B(_1643_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4634_ (.I(_0375_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4635_ (.A1(_0290_),
    .A2(_1644_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4636_ (.A1(_0281_),
    .A2(_0286_),
    .B(_0340_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4637_ (.A1(_0281_),
    .A2(_0286_),
    .B(_1646_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4638_ (.A1(_1645_),
    .A2(_1647_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4639_ (.A1(_0270_),
    .A2(_1644_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4640_ (.A1(_0288_),
    .A2(_0294_),
    .B(_0340_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4641_ (.A1(_0288_),
    .A2(_0294_),
    .B(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4642_ (.A1(_1648_),
    .A2(_1650_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4643_ (.A1(_0277_),
    .A2(_0296_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4644_ (.A1(_0277_),
    .A2(_0296_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4645_ (.A1(_1651_),
    .A2(_0347_),
    .A3(_1652_),
    .B1(_0397_),
    .B2(_0263_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4646_ (.A1(_0299_),
    .A2(_1651_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4647_ (.A1(_0297_),
    .A2(_0268_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4648_ (.A1(_1653_),
    .A2(_1654_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4649_ (.A1(_0254_),
    .A2(_1642_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4650_ (.A1(_0341_),
    .A2(_1655_),
    .B(_1656_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4651_ (.A1(_0261_),
    .A2(_0269_),
    .A3(_0301_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4652_ (.A1(_0269_),
    .A2(_0301_),
    .B(_0261_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4653_ (.A1(_1657_),
    .A2(_0347_),
    .A3(_1658_),
    .B1(_0397_),
    .B2(_0598_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4654_ (.A1(_0257_),
    .A2(_1657_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4655_ (.A1(_1659_),
    .A2(_0304_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4656_ (.A1(_0240_),
    .A2(_1642_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4657_ (.A1(_0341_),
    .A2(_1660_),
    .B(_1661_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4658_ (.A1(_0231_),
    .A2(_1644_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4659_ (.A1(_0306_),
    .A2(_0259_),
    .A3(_0330_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4660_ (.A1(_0308_),
    .A2(_1640_),
    .A3(_1663_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4661_ (.A1(_1662_),
    .A2(_1664_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4662_ (.A1(_0225_),
    .A2(_1644_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4663_ (.A1(_0244_),
    .A2(_0308_),
    .A3(_0310_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4664_ (.A1(_0332_),
    .A2(_1640_),
    .A3(_1666_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4665_ (.A1(_1665_),
    .A2(_1667_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4666_ (.A1(_0216_),
    .A2(_1642_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4667_ (.A1(_0235_),
    .A2(_0332_),
    .A3(_0333_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4668_ (.A1(_0313_),
    .A2(_1640_),
    .A3(_1669_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4669_ (.A1(_1668_),
    .A2(_1670_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4670_ (.A1(_0328_),
    .A2(_0334_),
    .A3(_0314_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4671_ (.I(_0213_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4672_ (.A1(_0316_),
    .A2(_0347_),
    .A3(_1671_),
    .B1(_0397_),
    .B2(_1672_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4673_ (.D(_0008_),
    .CLK(net89),
    .Q(\Control_Unit.T[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4674_ (.D(_0009_),
    .CLK(net89),
    .Q(\Control_Unit.T[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4675_ (.D(_0010_),
    .CLK(net90),
    .Q(\Control_Unit.T[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4676_ (.D(_0011_),
    .CLK(net92),
    .Q(\Control_Unit.T[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4677_ (.D(_0012_),
    .CLK(net92),
    .Q(\Control_Unit.T[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4678_ (.D(_0013_),
    .CLK(net110),
    .Q(\Control_Unit.T[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4679_ (.D(_0014_),
    .CLK(net110),
    .Q(\Control_Unit.T[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4680_ (.D(_0015_),
    .CLK(net110),
    .Q(\Control_Unit.T[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4681_ (.D(_0016_),
    .CLK(net111),
    .Q(\Control_Unit.T[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4682_ (.D(_0017_),
    .CLK(net115),
    .Q(\Control_Unit.T[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4683_ (.D(_0018_),
    .CLK(net111),
    .Q(\Control_Unit.T[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4684_ (.D(_0019_),
    .CLK(net98),
    .Q(\Control_Unit.T[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4685_ (.D(_0020_),
    .CLK(net98),
    .Q(\Control_Unit.T[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4686_ (.D(_0021_),
    .CLK(net106),
    .Q(\Control_Unit.T[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4687_ (.D(_0022_),
    .CLK(net105),
    .Q(\Control_Unit.T[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4688_ (.D(_0023_),
    .CLK(net97),
    .Q(\Control_Unit.T[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4689_ (.D(_0024_),
    .CLK(net96),
    .Q(\Control_Unit.T[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4690_ (.D(_0025_),
    .CLK(net85),
    .Q(\Control_Unit.T[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4691_ (.D(_0026_),
    .CLK(net96),
    .Q(\Control_Unit.T[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4692_ (.D(_0027_),
    .CLK(net99),
    .Q(\Control_Unit.T[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4693_ (.D(_0028_),
    .CLK(net52),
    .Q(\Control_Unit.cont[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4694_ (.D(_0029_),
    .CLK(net52),
    .Q(\Control_Unit.cont[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4695_ (.D(_0030_),
    .CLK(net52),
    .Q(\Control_Unit.cont[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4696_ (.D(_0031_),
    .CLK(net52),
    .Q(\Control_Unit.cont[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4697_ (.D(_0032_),
    .CLK(net54),
    .Q(\Control_Unit.cont[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4698_ (.D(_0033_),
    .CLK(net54),
    .Q(\Control_Unit.cont[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4699_ (.D(_0034_),
    .CLK(net59),
    .Q(\Control_Unit.cont[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4700_ (.D(_0035_),
    .CLK(net59),
    .Q(\Control_Unit.cont[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4701_ (.D(_0036_),
    .CLK(net57),
    .Q(\Control_Unit.cont[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4702_ (.D(_0037_),
    .CLK(net57),
    .Q(\Control_Unit.cont[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4703_ (.D(_0038_),
    .CLK(net57),
    .Q(\Control_Unit.cont[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4704_ (.D(_0039_),
    .CLK(net71),
    .Q(\Control_Unit.cont[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4705_ (.D(_0040_),
    .CLK(net58),
    .Q(\Control_Unit.cont[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4706_ (.D(_0041_),
    .CLK(net71),
    .Q(\Control_Unit.cont[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4707_ (.D(_0042_),
    .CLK(net74),
    .Q(\Control_Unit.cont[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4708_ (.D(_0043_),
    .CLK(net90),
    .Q(\Control_Unit.cont[15] ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _4709_ (.D(_0152_),
    .Q(\Control_Unit.Rc ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _4710_ (.D(_0002_),
    .Q(\Control_Unit.Rx ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _4711_ (.D(_0005_),
    .Q(\Control_Unit.Mc ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _4712_ (.D(_0003_),
    .Q(\Control_Unit.Mq ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _4713_ (.D(_0006_),
    .Q(\Control_Unit.Mt ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _4714_ (.D(_0001_),
    .Q(\Control_Unit.Mx ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _4715_ (.D(_0004_),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _4716_ (.D(_0000_),
    .Q(\Control_Unit.Rcont ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4717_ (.D(\Control_Unit.futuro[0] ),
    .CLK(net58),
    .Q(\Control_Unit.presente[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4718_ (.D(\Control_Unit.futuro[1] ),
    .CLK(net57),
    .Q(\Control_Unit.presente[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4719_ (.D(\Control_Unit.futuro[2] ),
    .CLK(net71),
    .Q(\Control_Unit.presente[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4720_ (.D(_0044_),
    .CLK(net77),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4721_ (.D(_0045_),
    .CLK(net77),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4722_ (.D(_0046_),
    .CLK(net67),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4723_ (.D(_0047_),
    .CLK(net67),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4724_ (.D(_0048_),
    .CLK(net77),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4725_ (.D(_0049_),
    .CLK(net78),
    .Q(net46));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4726_ (.D(_0050_),
    .CLK(net78),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4727_ (.D(_0051_),
    .CLK(net78),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4728_ (.D(_0052_),
    .CLK(net79),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4729_ (.D(_0053_),
    .CLK(net78),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4730_ (.D(_0054_),
    .CLK(net79),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4731_ (.D(_0055_),
    .CLK(net82),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4732_ (.D(_0056_),
    .CLK(net82),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4733_ (.D(_0057_),
    .CLK(net82),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4734_ (.D(_0058_),
    .CLK(net82),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4735_ (.D(_0059_),
    .CLK(net85),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4736_ (.D(_0060_),
    .CLK(net96),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4737_ (.D(_0061_),
    .CLK(net85),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4738_ (.D(_0062_),
    .CLK(net97),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4739_ (.D(_0063_),
    .CLK(net101),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4740_ (.D(_0064_),
    .CLK(net97),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4741_ (.D(_0065_),
    .CLK(net101),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4742_ (.D(_0066_),
    .CLK(net101),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4743_ (.D(_0067_),
    .CLK(net102),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4744_ (.D(_0068_),
    .CLK(net102),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4745_ (.D(_0069_),
    .CLK(net103),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4746_ (.D(_0070_),
    .CLK(net103),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4747_ (.D(_0071_),
    .CLK(net102),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4748_ (.D(_0072_),
    .CLK(net101),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4749_ (.D(_0073_),
    .CLK(net97),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4750_ (.D(_0074_),
    .CLK(net102),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4751_ (.D(_0075_),
    .CLK(net96),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4752_ (.D(_0076_),
    .CLK(net77),
    .Q(\Control_Unit.Q[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4753_ (.D(_0077_),
    .CLK(net55),
    .Q(\Control_Unit.Q[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4754_ (.D(_0078_),
    .CLK(net53),
    .Q(\Control_Unit.Q[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4755_ (.D(_0079_),
    .CLK(net53),
    .Q(\Control_Unit.Q[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4756_ (.D(_0080_),
    .CLK(net80),
    .Q(\Control_Unit.Q[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4757_ (.D(_0081_),
    .CLK(net53),
    .Q(\Control_Unit.Q[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4758_ (.D(_0082_),
    .CLK(net55),
    .Q(\Control_Unit.Q[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4759_ (.D(_0083_),
    .CLK(net55),
    .Q(\Control_Unit.Q[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4760_ (.D(_0084_),
    .CLK(net56),
    .Q(\Control_Unit.Q[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4761_ (.D(_0085_),
    .CLK(net56),
    .Q(\Control_Unit.Q[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4762_ (.D(_0086_),
    .CLK(net71),
    .Q(\Control_Unit.Q[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4763_ (.D(_0087_),
    .CLK(net72),
    .Q(\Control_Unit.Q[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4764_ (.D(_0088_),
    .CLK(net72),
    .Q(\Control_Unit.Q[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4765_ (.D(_0089_),
    .CLK(net73),
    .Q(\Control_Unit.Q[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4766_ (.D(_0090_),
    .CLK(net73),
    .Q(\Control_Unit.Q[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4767_ (.D(_0091_),
    .CLK(net90),
    .Q(\Control_Unit.Q[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4768_ (.D(_0092_),
    .CLK(net91),
    .Q(\Control_Unit.Q[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4769_ (.D(_0093_),
    .CLK(net93),
    .Q(\Control_Unit.Q[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4770_ (.D(_0094_),
    .CLK(net112),
    .Q(\Control_Unit.Q[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4771_ (.D(_0095_),
    .CLK(net112),
    .Q(\Control_Unit.Q[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4772_ (.D(_0096_),
    .CLK(net114),
    .Q(\Control_Unit.Q[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4773_ (.D(_0097_),
    .CLK(net114),
    .Q(\Control_Unit.Q[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4774_ (.D(_0098_),
    .CLK(net114),
    .Q(\Control_Unit.Q[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4775_ (.D(_0099_),
    .CLK(net106),
    .Q(\Control_Unit.Q[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4776_ (.D(_0100_),
    .CLK(net107),
    .Q(\Control_Unit.Q[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4777_ (.D(_0101_),
    .CLK(net107),
    .Q(\Control_Unit.Q[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4778_ (.D(_0102_),
    .CLK(net107),
    .Q(\Control_Unit.Q[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4779_ (.D(_0103_),
    .CLK(net106),
    .Q(\Control_Unit.Q[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4780_ (.D(_0104_),
    .CLK(net83),
    .Q(\Control_Unit.Q[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4781_ (.D(_0105_),
    .CLK(net83),
    .Q(\Control_Unit.Q[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4782_ (.D(_0106_),
    .CLK(net86),
    .Q(\Control_Unit.Q[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4783_ (.D(_0107_),
    .CLK(net87),
    .Q(\Control_Unit.Q[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4784_ (.D(_0108_),
    .CLK(net67),
    .Q(\Control_Unit.C[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4785_ (.D(_0109_),
    .CLK(net61),
    .Q(\Control_Unit.C[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4786_ (.D(_0110_),
    .CLK(net62),
    .Q(\Control_Unit.C[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4787_ (.D(_0111_),
    .CLK(net61),
    .Q(\Control_Unit.C[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4788_ (.D(_0112_),
    .CLK(net62),
    .Q(\Control_Unit.C[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4789_ (.D(_0113_),
    .CLK(net63),
    .Q(\Control_Unit.C[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4790_ (.D(_0114_),
    .CLK(net63),
    .Q(\Control_Unit.C[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4791_ (.D(_0115_),
    .CLK(net63),
    .Q(\Control_Unit.C[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4792_ (.D(_0116_),
    .CLK(net63),
    .Q(\Control_Unit.C[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4793_ (.D(_0117_),
    .CLK(net64),
    .Q(\Control_Unit.C[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4794_ (.D(_0118_),
    .CLK(net72),
    .Q(\Control_Unit.C[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4795_ (.D(_0119_),
    .CLK(net72),
    .Q(\Control_Unit.C[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4796_ (.D(_0120_),
    .CLK(net73),
    .Q(\Control_Unit.C[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4797_ (.D(_0121_),
    .CLK(net89),
    .Q(\Control_Unit.C[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4798_ (.D(_0122_),
    .CLK(net91),
    .Q(\Control_Unit.C[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4799_ (.D(_0123_),
    .CLK(net92),
    .Q(\Control_Unit.C[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4800_ (.D(_0124_),
    .CLK(net92),
    .Q(\Control_Unit.C[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4801_ (.D(_0125_),
    .CLK(net93),
    .Q(\Control_Unit.C[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4802_ (.D(_0126_),
    .CLK(net113),
    .Q(\Control_Unit.C[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4803_ (.D(_0127_),
    .CLK(net113),
    .Q(\Control_Unit.C[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4804_ (.D(_0128_),
    .CLK(net110),
    .Q(\Control_Unit.C[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4805_ (.D(_0129_),
    .CLK(net114),
    .Q(\Control_Unit.C[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4806_ (.D(_0130_),
    .CLK(net99),
    .Q(\Control_Unit.C[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4807_ (.D(_0131_),
    .CLK(net100),
    .Q(\Control_Unit.C[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4808_ (.D(_0132_),
    .CLK(net98),
    .Q(\Control_Unit.C[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4809_ (.D(_0133_),
    .CLK(net106),
    .Q(\Control_Unit.C[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4810_ (.D(_0134_),
    .CLK(net98),
    .Q(\Control_Unit.C[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4811_ (.D(_0135_),
    .CLK(net99),
    .Q(\Control_Unit.C[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4812_ (.D(_0136_),
    .CLK(net84),
    .Q(\Control_Unit.C[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4813_ (.D(_0137_),
    .CLK(net85),
    .Q(\Control_Unit.C[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4814_ (.D(_0138_),
    .CLK(net84),
    .Q(\Control_Unit.C[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4815_ (.D(_0139_),
    .CLK(net87),
    .Q(\Control_Unit.C[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4816_ (.D(_0140_),
    .CLK(net68),
    .Q(\Control_Unit.T[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4817_ (.D(_0141_),
    .CLK(net67),
    .Q(\Control_Unit.T[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4818_ (.D(_0142_),
    .CLK(net61),
    .Q(\Control_Unit.T[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4819_ (.D(_0143_),
    .CLK(net61),
    .Q(\Control_Unit.T[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4820_ (.D(_0144_),
    .CLK(net68),
    .Q(\Control_Unit.T[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4821_ (.D(_0145_),
    .CLK(net68),
    .Q(\Control_Unit.T[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4822_ (.D(_0146_),
    .CLK(net69),
    .Q(\Control_Unit.T[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4823_ (.D(_0147_),
    .CLK(net81),
    .Q(\Control_Unit.T[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4824_ (.D(_0148_),
    .CLK(net64),
    .Q(\Control_Unit.T[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4825_ (.D(_0149_),
    .CLK(net69),
    .Q(\Control_Unit.T[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4826_ (.D(_0150_),
    .CLK(net81),
    .Q(\Control_Unit.T[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4827_ (.D(_0151_),
    .CLK(net89),
    .Q(\Control_Unit.T[11] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(clk),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input2 (.I(n[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(n[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(n[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(n[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(n[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input7 (.I(n[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input8 (.I(n[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(n[1]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(n[2]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input11 (.I(n[3]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(n[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(n[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(n[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(n[7]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(n[8]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input17 (.I(n[9]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(start),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(X[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(X[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(X[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(X[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(X[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(X[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(X[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(X[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(X[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(X[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(X[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(X[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(X[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(X[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(X[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(X[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(X[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(X[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(X[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(X[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(X[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(X[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(X[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(X[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(X[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(X[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(X[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output46 (.I(net46),
    .Z(X[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output47 (.I(net47),
    .Z(X[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output48 (.I(net48),
    .Z(X[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output49 (.I(net49),
    .Z(X[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output50 (.I(net50),
    .Z(X[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output51 (.I(net51),
    .Z(b));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout52 (.I(net54),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout53 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout54 (.I(net55),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout55 (.I(net60),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout56 (.I(net60),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout57 (.I(net58),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout58 (.I(net59),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout59 (.I(net60),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net76),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout61 (.I(net66),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout62 (.I(net66),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout63 (.I(net65),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout65 (.I(net66),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net70),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout67 (.I(net69),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout68 (.I(net69),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout69 (.I(net70),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout70 (.I(net75),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout71 (.I(net74),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout72 (.I(net73),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout73 (.I(net74),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net76),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout76 (.I(net119),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout77 (.I(net80),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout78 (.I(net80),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout79 (.I(net80),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout80 (.I(net81),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout81 (.I(net88),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout82 (.I(net84),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout84 (.I(net86),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout85 (.I(net86),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout86 (.I(net87),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout88 (.I(net95),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout89 (.I(net90),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout90 (.I(net94),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout91 (.I(net94),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout92 (.I(net93),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net94),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout94 (.I(net95),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout95 (.I(net118),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout96 (.I(net100),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout97 (.I(net100),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout98 (.I(net99),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout99 (.I(net100),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout100 (.I(net109),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout101 (.I(net105),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout102 (.I(net104),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout103 (.I(net104),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout104 (.I(net105),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout105 (.I(net108),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout106 (.I(net107),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout107 (.I(net108),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout108 (.I(net109),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout109 (.I(net117),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout110 (.I(net112),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout111 (.I(net112),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout112 (.I(net116),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net116),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout114 (.I(net115),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout115 (.I(net116),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout116 (.I(net117),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout117 (.I(net118),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout118 (.I(net119),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout119 (.I(net1),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(\Control_Unit.C[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A2 (.I(\Control_Unit.C[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A2 (.I(\Control_Unit.C[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__I (.I(\Control_Unit.C[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A2 (.I(\Control_Unit.C[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A2 (.I(\Control_Unit.C[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__I (.I(\Control_Unit.C[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A2 (.I(\Control_Unit.C[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(\Control_Unit.C[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A2 (.I(\Control_Unit.C[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__I (.I(\Control_Unit.C[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A2 (.I(\Control_Unit.C[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A2 (.I(\Control_Unit.C[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A2 (.I(\Control_Unit.C[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__I (.I(\Control_Unit.C[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A2 (.I(\Control_Unit.C[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A2 (.I(\Control_Unit.C[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__I (.I(\Control_Unit.C[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A2 (.I(\Control_Unit.C[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A2 (.I(\Control_Unit.C[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A2 (.I(\Control_Unit.C[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__I (.I(\Control_Unit.C[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A2 (.I(\Control_Unit.C[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A2 (.I(\Control_Unit.C[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A2 (.I(\Control_Unit.C[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__I (.I(\Control_Unit.C[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A2 (.I(\Control_Unit.C[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A2 (.I(\Control_Unit.C[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A2 (.I(\Control_Unit.C[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__I (.I(\Control_Unit.C[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A2 (.I(\Control_Unit.C[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A2 (.I(\Control_Unit.C[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__I (.I(\Control_Unit.C[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(\Control_Unit.C[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(\Control_Unit.C[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__I (.I(\Control_Unit.C[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__I (.I(\Control_Unit.C[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A2 (.I(\Control_Unit.C[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A2 (.I(\Control_Unit.C[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A2 (.I(\Control_Unit.C[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__I (.I(\Control_Unit.C[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__B (.I(\Control_Unit.C[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(\Control_Unit.C[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A2 (.I(\Control_Unit.C[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A3 (.I(\Control_Unit.C[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(\Control_Unit.C[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A2 (.I(\Control_Unit.C[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A1 (.I(\Control_Unit.C[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__I (.I(\Control_Unit.C[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A2 (.I(\Control_Unit.C[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__I (.I(\Control_Unit.C[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A2 (.I(\Control_Unit.C[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A2 (.I(\Control_Unit.C[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__I (.I(\Control_Unit.C[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A2 (.I(\Control_Unit.C[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(\Control_Unit.C[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A2 (.I(\Control_Unit.C[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__I (.I(\Control_Unit.C[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(\Control_Unit.C[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A2 (.I(\Control_Unit.C[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A2 (.I(\Control_Unit.C[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__I (.I(\Control_Unit.C[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(\Control_Unit.C[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A2 (.I(\Control_Unit.C[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A2 (.I(\Control_Unit.C[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__I (.I(\Control_Unit.C[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__I (.I(\Control_Unit.Mq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__I (.I(\Control_Unit.Mq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A2 (.I(\Control_Unit.Mq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__I (.I(\Control_Unit.Mq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__I (.I(\Control_Unit.Mx ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A2 (.I(\Control_Unit.Mx ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__I (.I(\Control_Unit.Mx ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__I (.I(\Control_Unit.Q[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(\Control_Unit.Q[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A1 (.I(\Control_Unit.Q[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A3 (.I(\Control_Unit.Q[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(\Control_Unit.Q[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__I (.I(\Control_Unit.Q[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A1 (.I(\Control_Unit.Q[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A3 (.I(\Control_Unit.Q[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__I (.I(\Control_Unit.Q[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A2 (.I(\Control_Unit.Q[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(\Control_Unit.Q[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__A3 (.I(\Control_Unit.Q[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A2 (.I(\Control_Unit.Q[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__I (.I(\Control_Unit.Q[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(\Control_Unit.Q[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A3 (.I(\Control_Unit.Q[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A2 (.I(\Control_Unit.Q[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__I (.I(\Control_Unit.Q[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A1 (.I(\Control_Unit.Q[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A3 (.I(\Control_Unit.Q[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__I (.I(\Control_Unit.Q[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A2 (.I(\Control_Unit.Q[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A1 (.I(\Control_Unit.Q[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A3 (.I(\Control_Unit.Q[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A2 (.I(\Control_Unit.Q[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__I (.I(\Control_Unit.Q[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A2 (.I(\Control_Unit.Q[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A1 (.I(\Control_Unit.Q[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__I (.I(\Control_Unit.Q[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A1 (.I(\Control_Unit.Q[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A3 (.I(\Control_Unit.Q[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__I (.I(\Control_Unit.Q[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A3 (.I(\Control_Unit.Q[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A1 (.I(\Control_Unit.Q[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A3 (.I(\Control_Unit.Q[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__I (.I(\Control_Unit.Q[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A1 (.I(\Control_Unit.Q[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A3 (.I(\Control_Unit.Q[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(\Control_Unit.Q[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__I (.I(\Control_Unit.Q[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A1 (.I(\Control_Unit.Q[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A3 (.I(\Control_Unit.Q[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A2 (.I(\Control_Unit.Q[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A2 (.I(\Control_Unit.Q[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__I (.I(\Control_Unit.Q[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A3 (.I(\Control_Unit.Q[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A2 (.I(\Control_Unit.Q[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__I (.I(\Control_Unit.Q[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__A1 (.I(\Control_Unit.Q[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A3 (.I(\Control_Unit.Q[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(\Control_Unit.Q[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__I (.I(\Control_Unit.Q[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A1 (.I(\Control_Unit.Q[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A3 (.I(\Control_Unit.Q[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(\Control_Unit.Rc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__I (.I(\Control_Unit.Rc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__A1 (.I(\Control_Unit.Rc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__I (.I(\Control_Unit.Rc ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__A1 (.I(\Control_Unit.Rcont ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__I (.I(\Control_Unit.Rcont ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__I (.I(\Control_Unit.Rcont ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__I (.I(\Control_Unit.T[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A2 (.I(\Control_Unit.T[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A2 (.I(\Control_Unit.T[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A2 (.I(\Control_Unit.T[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A3 (.I(\Control_Unit.T[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__I (.I(\Control_Unit.T[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A3 (.I(\Control_Unit.T[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A1 (.I(\Control_Unit.T[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__I (.I(\Control_Unit.T[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__A1 (.I(\Control_Unit.T[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A1 (.I(\Control_Unit.T[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(\Control_Unit.T[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A2 (.I(\Control_Unit.T[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__I (.I(\Control_Unit.T[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A1 (.I(\Control_Unit.T[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A1 (.I(\Control_Unit.T[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__A2 (.I(\Control_Unit.T[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__I (.I(\Control_Unit.T[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(\Control_Unit.cont[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A1 (.I(\Control_Unit.cont[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__I (.I(\Control_Unit.cont[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__I (.I(\Control_Unit.cont[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(\Control_Unit.cont[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__I (.I(\Control_Unit.cont[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__I (.I(\Control_Unit.cont[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A1 (.I(\Control_Unit.cont[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__I (.I(\Control_Unit.cont[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__I (.I(\Control_Unit.cont[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A1 (.I(\Control_Unit.cont[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__I (.I(\Control_Unit.cont[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A2 (.I(\Control_Unit.cont[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__I (.I(\Control_Unit.cont[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__I (.I(\Control_Unit.cont[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A1 (.I(\Control_Unit.cont[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__I (.I(\Control_Unit.cont[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A1 (.I(\Control_Unit.cont[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__I (.I(\Control_Unit.cont[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__D (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__D (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__D (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__D (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__D (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__D (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__D (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__D (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__D (.I(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__D (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__D (.I(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__D (.I(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__D (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__D (.I(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__D (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__D (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__D (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__B (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__A2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__B2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__A2 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__B (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__B1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__A2 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__A2 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__I (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A2 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A2 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A2 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__A2 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A2 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__A2 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__A3 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__A2 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__A2 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A1 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A1 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__A1 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__I (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A2 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A2 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__I (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__A2 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__B (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__A3 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__A3 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__B (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__B (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__B (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__I (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__B1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__A3 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__B (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__B (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__B (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__B (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__B1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__B1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__C (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__B (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__I (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__I (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__A3 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__B1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__I (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__I (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A3 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__B (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__B (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__I (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__I (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__A3 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__B1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__B1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__B1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__B1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A3 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__A2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__B (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__A2 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__A2 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__B2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__C (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__B (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__B (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__S (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__I (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__B (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__B (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__B (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__S (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__I (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__B2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__B2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__B2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__B (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__I (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__I (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__I (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__I (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__I (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__I (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__I (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__B1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__B1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__B1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__B1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__B (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A3 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A3 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__B (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__B (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__B (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A3 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__I (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__B1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__B (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__B (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__A2 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A2 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A2 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__B2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A3 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__B (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A3 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A3 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__B1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__B1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__B1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__B1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__B (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__B (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__B (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__B (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__B (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__B2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__B (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__B2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A3 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__I (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__B (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__B1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__B1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__B1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__B1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__B2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A3 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__B (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__B2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__B (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__B (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__B (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__B (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__B (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__B2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A4 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__B (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__B2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__I (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__B (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__B1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__B1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__B1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__S (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__B2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__B1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__I (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__I (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__I (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__B1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__B1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__B (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__I (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__I (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A2 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A2 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A3 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A3 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__B (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__B (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__B2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__B (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__B1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__B1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__B1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__I (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A3 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A3 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__I (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__I (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__B1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__B1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__B (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__B1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__B2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__I (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A2 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A2 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__C (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__B (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A3 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__B (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__B (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__I (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A3 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A2 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A3 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__I (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__I (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__B (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__B (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__I (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__I (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A2 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A2 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__B (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__B (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__B1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__B1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__B1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A3 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__B (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__B (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__B (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__B1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__B1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__I (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__B (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__B (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__I (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__B (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__B1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__B1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A3 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A3 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A4 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__I (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A3 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A2 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__B (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__A2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__B1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__B2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__A2 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A2 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__B2 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__I (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__B2 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__B2 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A4 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__B2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__B2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__B2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A1 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A1 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A3 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__B2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A4 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__B2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A4 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A3 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__I (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__A3 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__B (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__C (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__A1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__I (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__I (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__I (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__I (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__I (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__I (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__I (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__I (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__I (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A1 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A1 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__I (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__I (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__I (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__I (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__I (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A1 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__I (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A3 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__I (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__I1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A3 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A3 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__I (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A2 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A2 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A2 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A3 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__I (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__I (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__I (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A1 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A1 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__I (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A2 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__I (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__B (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A1 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__B (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__B (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A1 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__I (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A2 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__I (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__I0 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__I (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__I1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__I (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A1 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A1 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__I (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A3 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__I (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__I (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__I (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__B (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__A1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__B (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A1 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A3 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A2 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__I0 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__I (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__B (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__B (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A3 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__I (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__I (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__I (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A3 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__I (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__B1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__I (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__A3 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A1 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A3 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__I (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__A1 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__I (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A3 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A3 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__B2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__I (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A1 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__I (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__I (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__I (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__I (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__B2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__I (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A1 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__I (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__I (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__I1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A1 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__A2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A4 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__I (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__I (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__I (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__I (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__I (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__I (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__B (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A2 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A1 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__A1 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__C (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A1 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A1 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A1 (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A2 (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A1 (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__I0 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__I (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A2 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__S (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__I (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__I (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A1 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A1 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__I (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__A3 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__I (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__B1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__A1 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A1 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__I1 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A2 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__B1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A2 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A2 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__B1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__B1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A1 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__I (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A1 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__I1 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__B1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__A1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__I0 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__I (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__A2 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__A1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__I1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__B2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3027__B2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__B (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__I (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A1 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A1 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A1 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__I (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__A1 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__A1 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A1 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A1 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__I (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__A1 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__B2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__I (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__A1 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__A2 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A1 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A1 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__A2 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A2 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__B2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__B1 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__B1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A2 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__I (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__B2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A3 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__I (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__I (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__A2 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A2 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A2 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A1 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__I (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__C (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A2 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__A2 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__I (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__A3 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A2 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__A4 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__I (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A1 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__I (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__I (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__I (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__I (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A2 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A2 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__I (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A3 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A2 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__I (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A3 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A1 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A4 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A3 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A3 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__I (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A2 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__I (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__I (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A2 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__A2 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A4 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A1 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__I (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A1 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A1 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A3 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A4 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A2 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__I (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A2 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A2 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A3 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A3 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A4 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__I (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__I (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__B2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__I (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__I (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A3 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__I (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A1 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A1 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__I (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__I (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__I (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A1 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__A3 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__I (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__C (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__I (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__I (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A2 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__B2 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A2 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A2 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A1 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__I (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__A1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A2 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A2 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A2 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__B2 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__I (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__I (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A2 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A1 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__A1 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A1 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__A2 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A2 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__B1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__B (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__A2 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__B (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__C (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__A3 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__B1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__B2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A2 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A2 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A3 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__I (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__A2 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A2 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__I (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__A1 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__I (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__I (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__B (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__B2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__I (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__A3 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A3 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A4 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A1 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__I (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__A1 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__A3 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A3 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__B (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__A3 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A2 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A2 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__A1 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A3 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A1 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__A1 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__A1 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__A2 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__B (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A2 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__A3 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__B (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__B (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A2 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A2 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__C (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A2 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A1 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__A1 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3027__A1 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A1 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A3 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__B1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(n[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(n[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(n[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(n[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(n[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(n[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(n[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(n[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(n[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(n[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(n[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(n[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(n[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(n[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(n[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(n[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(start));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__B1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__B2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__B2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A3 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__B2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__B2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__B2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__B2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__CLK (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__CLK (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__CLK (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout61_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout77_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout80_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__CLK (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__CLK (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__CLK (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__CLK (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__CLK (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__CLK (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout114_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout76_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
endmodule

