* NGSPICE file created from suma_mult_TOP.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_1 D E RN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

.subckt suma_mult_TOP X[0] X[10] X[11] X[12] X[13] X[14] X[15] X[16] X[17] X[18] X[19]
+ X[1] X[20] X[21] X[22] X[23] X[24] X[25] X[26] X[27] X[28] X[29] X[2] X[30] X[31]
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] b clk n[0] n[10] n[11] n[12] n[13] n[14] n[15]
+ n[1] n[2] n[3] n[4] n[5] n[6] n[7] n[8] n[9] start vdd vss
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3140__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3155_ _0274_ _0275_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout56_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3086_ _2111_ Control_Unit.T\[9\] _2050_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3988_ _1033_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2939_ _2265_ _2243_ _2266_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_10_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2954__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4609_ _0490_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4459__A1 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3131__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2863__I _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2642__B1 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3673__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A1 Control_Unit.C\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ _1803_ _0557_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3842_ Control_Unit.Q\[29\] _0918_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3773_ _0839_ _0845_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2936__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2724_ _2049_ _2052_ _2048_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2655_ Control_Unit.C\[23\] _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4325_ _1358_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2586_ _1914_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3361__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout116 net117 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout105 net108 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ _1172_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4187_ _1242_ _1244_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3207_ _0319_ _0349_ _1881_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3138_ _1801_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3069_ Control_Unit.T\[11\] _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3104__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2918__A1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2394__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3591__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout106_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2440_ Control_Unit.cont\[3\] _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2371_ net5 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4110_ _1171_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4041_ _2055_ _1105_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3548__B _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3825_ _0492_ _1996_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3756_ _0464_ Control_Unit.C\[24\] Control_Unit.Q\[24\] _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ _1868_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3687_ _0522_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2638_ _1966_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2678__I _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3334__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2569_ _1764_ _1850_ _1854_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2688__A3 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ Control_Unit.Mc _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4239_ _0814_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3325__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4289__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3628__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3610_ _0696_ _0702_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4590_ _1353_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ Control_Unit.T\[9\] _2000_ Control_Unit.Q\[9\] _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_7_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3564__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3316__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3472_ _2015_ _0270_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2423_ _1714_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2354_ _1684_ _0007_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3867__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4024_ _1067_ _1069_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3278__B _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3808_ _0865_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4788_ _0112_ net62 Control_Unit.C\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3739_ _0457_ Control_Unit.C\[22\] _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3086__A3 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__A2 Control_Unit.Q\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3546__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3849__A2 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2521__A2 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2972_ _2294_ _2298_ _2299_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4711_ _0005_ _4711_/E _4711_/RN Control_Unit.Mc vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__2588__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _1648_ _1650_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4573_ _1422_ _1593_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3524_ net49 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3455_ _2016_ _0290_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2406_ Control_Unit.cont\[13\] _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3386_ _0508_ _2145_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout86_I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2337_ _1673_ _1674_ Control_Unit.presente\[0\] _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3068__A3 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4007_ Control_Unit.Q\[9\] _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4265__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2691__I Control_Unit.C\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3776__A1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3059__A3 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4784__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4192__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3240_ _0367_ _0370_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3171_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4247__A2 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _2282_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2886_ _1861_ _1864_ _1869_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4625_ _0941_ _0532_ _0340_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4556_ _1578_ _1579_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2733__A2 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3507_ _0604_ _0608_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4487_ _1506_ _1511_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3438_ Control_Unit.Q\[1\] _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3291__B _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3369_ _0492_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2686__I Control_Unit.C\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3997__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput42 net42 X[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput31 net31 X[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput20 net20 X[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4252__S _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2740_ _2067_ _2068_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2963__A2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2671_ Control_Unit.C\[9\] _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3376__B _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4410_ _1766_ _1430_ _1445_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3912__A1 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4341_ _1372_ _1381_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _1306_ _1317_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3223_ _0348_ _0337_ _0355_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3140__A2 Control_Unit.T\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3154_ _0297_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3085_ _0223_ _0228_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2651__A1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3987_ Control_Unit.Q\[8\] _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2403__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2938_ _2241_ _2242_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2954__A2 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4156__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2869_ _2190_ _2193_ _2196_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4608_ _1620_ _1623_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4539_ _1992_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2642__B2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4822__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3122__A2 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2881__A1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4046__I _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4622__A2 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2633__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3910_ _0971_ _0980_ _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3841_ Control_Unit.T\[29\] _1995_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3772_ _0840_ _0844_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4386__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2723_ _2050_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2654_ Control_Unit.C\[20\] _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2585_ _1769_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4324_ Control_Unit.C\[2\] _1795_ _1803_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout117 net118 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout106 net107 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4255_ _1174_ _1171_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4186_ _1242_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3206_ Control_Unit.T\[13\] _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2872__A1 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3137_ _1814_ _0278_ _0280_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3068_ _1681_ _1679_ _2185_ _0212_ Control_Unit.futuro\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_35_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2624__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__B1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A1 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4129__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3104__A2 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2615__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2394__A3 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2370_ _1695_ _1696_ _1697_ _1698_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4040_ _1079_ _1085_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2854__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2606__A1 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4359__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3824_ _0492_ Control_Unit.C\[28\] _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3755_ _0835_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3031__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2706_ _2034_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3686_ _0773_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2637_ _1708_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2568_ _1866_ _1893_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2688__A4 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4307_ _0525_ _0941_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2499_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4238_ _1708_ _0768_ _0788_ _0797_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__3098__A1 _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4169_ _1213_ _1210_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4598__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3573__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3325__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3089__A1 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3540_ net50 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3471_ Control_Unit.T\[4\] _2008_ Control_Unit.Q\[4\] _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2422_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3316__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2353_ _1686_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4690__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4023_ _1087_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2827__B2 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2827__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4044__A3 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3807_ _0873_ _0880_ _0881_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4787_ _0111_ net61 Control_Unit.C\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3738_ _0457_ Control_Unit.C\[22\] _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3669_ _0427_ Control_Unit.C\[18\] Control_Unit.Q\[18\] _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4504__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2818__A1 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3491__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3794__A2 Control_Unit.C\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2754__B1 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2599__I _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2809__A1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3482__A1 Control_Unit.T\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2971_ _2056_ _2226_ _2236_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__3234__A1 Control_Unit.Rc vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4710_ _0002_ _4710_/E _4710_/RN Control_Unit.Rx vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _0288_ _0294_ _1649_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4572_ _1584_ _1436_ _1591_ _1595_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3523_ _0528_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3454_ _0557_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ Control_Unit.cont\[14\] _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3385_ _0506_ _0508_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2336_ Control_Unit.presente\[1\] _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_fanout79_I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4006_ _1055_ _0937_ _1056_ _1073_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3473__A1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3225__A1 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3528__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3662__B _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3170_ _0214_ _0219_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4049__I Control_Unit.Q\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3455__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3758__A2 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2954_ _2063_ _2280_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2885_ _1758_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _1634_ _1635_ _1636_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4183__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4555_ _1575_ _1576_ _1578_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3506_ _0570_ _0579_ _0605_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _1503_ _1462_ _1513_ _1516_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3437_ _0541_ _0542_ Control_Unit.T\[2\] _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3368_ Control_Unit.T\[29\] _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3299_ _0434_ _0429_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input11_I n[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3747__B _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput32 net32 X[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput43 net43 X[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput21 net21 X[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_49_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3685__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2488__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2670_ _1986_ _1994_ _1998_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4165__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3912__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4340_ _1371_ _1378_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4271_ Control_Unit.Q\[25\] _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3222_ _0350_ _0354_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I n[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3153_ _0266_ _0267_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3084_ _0224_ _0226_ _0227_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3428__A1 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3411__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2651__A2 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3986_ _0996_ _1053_ _1054_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2403__A2 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2937_ _1828_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2954__A3 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2868_ _1732_ _1873_ _2195_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_11_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4607_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2799_ _2072_ _2078_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4538_ _1557_ _1564_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4774__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2697__I _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4469_ _1498_ _1499_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3419__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4083__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3840_ Control_Unit.T\[29\] _1995_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3771_ _0850_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2397__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2722_ _1781_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3594__B1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4797__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2653_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3897__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2584_ _1828_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ _1357_ _1362_ _1363_ _1365_ _1360_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout118 net119 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout107 net108 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4254_ Control_Unit.Q\[24\] _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4185_ _1728_ _1221_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3205_ _0321_ _0325_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3136_ _1925_ _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout61_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3067_ _1973_ _0211_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3821__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3969_ _1020_ _1022_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4301__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4065__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2615__A2 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3879__A1 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4056__A1 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2606__A2 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3823_ _0495_ Control_Unit.C\[29\] Control_Unit.Q\[29\] _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4359__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3754_ _0836_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _1873_ _2030_ _2031_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3685_ _0754_ _0757_ _0763_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2636_ net8 _1887_ _1960_ _1963_ _1961_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2790__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2567_ _1894_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2498_ _1819_ _1815_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4306_ _1349_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4237_ _1291_ _1287_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3098__A2 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4168_ _1225_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4099_ _1144_ _1146_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3119_ _0262_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2533__A1 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3325__A3 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4038__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2834__B _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3261__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout111_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3470_ net45 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2421_ _1749_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2524__A1 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2352_ _1673_ _1685_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4022_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3252__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3806_ net39 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4786_ _0110_ net62 Control_Unit.C\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3737_ Control_Unit.Q\[22\] _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3668_ _0754_ _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3599_ Control_Unit.Q\[12\] _0692_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2619_ _1941_ _1946_ _1947_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4268__A1 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2818__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4708__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4440__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2754__B2 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4259__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2809__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3482__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2970_ _2295_ _2296_ _2297_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3234__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ _0288_ _0294_ _0340_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4571_ _1584_ _1594_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2745__A1 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3522_ _0582_ _0610_ _0622_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3453_ Control_Unit.C\[3\] Control_Unit.T\[3\] _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2404_ _1732_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3384_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2335_ Control_Unit.presente\[2\] _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4005_ _1070_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3473__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3225__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4769_ _0093_ net93 Control_Unit.Q\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2736__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4489__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4583__C _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4680__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3924__B1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3207__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2953_ _1763_ _1779_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2884_ _2209_ _2210_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3409__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ _1514_ _1633_ Control_Unit.C\[31\] _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4554_ _1990_ _1577_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3391__A1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3505_ _0593_ _0606_ _0591_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout91_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4485_ _1514_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3436_ Control_Unit.Q\[2\] _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3367_ _0486_ _0489_ _0494_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4238__A4 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3298_ Control_Unit.T\[19\] _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2957__A1 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2709__A1 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput33 net33 X[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput22 net22 X[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput44 net44 X[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3685__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3437__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2948__A1 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3373__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _1321_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3221_ _0343_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3152_ _0288_ _0294_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3083_ _2112_ _0225_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4625__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2636__B1 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2939__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3985_ _0611_ _1014_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3600__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ _2254_ _2258_ _2263_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2867_ _1890_ _2029_ _2194_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4606_ _1607_ _1606_ _1604_ _1621_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2798_ _2082_ _1913_ _2071_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4537_ _1558_ _1562_ _1563_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4468_ _1496_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3419_ _0525_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4399_ _1350_ _1434_ _1435_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3658__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4755__D _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3770_ Control_Unit.Q\[24\] _0851_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2721_ _1852_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3594__B2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3594__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2652_ Control_Unit.C\[21\] _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2583_ _1823_ _1911_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4322_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout119 net1 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4253_ _1305_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3204_ _0346_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4184_ _1218_ _1220_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3422__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3135_ _1812_ Control_Unit.T\[1\] _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3066_ _1676_ _2024_ _1673_ _1677_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_fanout54_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3282__B1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3578__B _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3297__C _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3968_ _0239_ _1024_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2919_ _2240_ _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3899_ _0953_ _0954_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4428__I _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3879__A2 Control_Unit.Q\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3242__I _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3500__A1 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4764__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3822_ net40 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3753_ _0821_ _0825_ _0828_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2704_ _2031_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3684_ _0759_ _0762_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2635_ net7 _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2790__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3417__I _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2566_ _1856_ _1860_ _1869_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4305_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2497_ _1825_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4236_ _1283_ _1285_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ _0383_ _1208_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4295__A2 Control_Unit.Q\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3118_ Control_Unit.T\[4\] _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4098_ _1144_ _1146_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3049_ _1964_ _2314_ _0192_ _0194_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_24_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__A2 _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3730__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4286__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4038__A2 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2406__I Control_Unit.cont\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout90 net94 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_31_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2420_ _1748_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout104_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2351_ _1677_ _1683_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2524__A2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4021_ _1075_ _1076_ _1086_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4785_ _0109_ net61 Control_Unit.C\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3805_ _0540_ _0883_ _0884_ _0885_ _0519_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3736_ _0456_ Control_Unit.C\[23\] Control_Unit.Q\[23\] _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_14_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3667_ _0744_ _0747_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3598_ _0318_ _2019_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2618_ _1691_ _1908_ _1945_ net13 _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2549_ _1874_ _1877_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4219_ _0940_ _1273_ _1275_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3057__I _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3219__B1 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3482__A3 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4570_ _0421_ _1593_ _1364_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2745__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3521_ _0617_ _0620_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3452_ Control_Unit.Q\[3\] _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2403_ _1708_ _1727_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3383_ Control_Unit.Rcont _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4004_ _1049_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3225__A3 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2433__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4768_ _0092_ net91 Control_Unit.Q\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4699_ _0034_ net59 Control_Unit.cont\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2736__A2 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3719_ _0765_ _0795_ _0805_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3933__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4489__A2 Control_Unit.C\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4825__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2424__A1 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2975__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3924__B2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4758__D _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__A1 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3207__A3 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2415__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2952_ _1766_ _1779_ _1782_ _2063_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2883_ _2209_ _2210_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4622_ Control_Unit.C\[31\] _1406_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4553_ _1991_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3915__A1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4484_ _1505_ _1501_ _1512_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3504_ _0585_ _0589_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3435_ Control_Unit.C\[2\] _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3425__I _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3366_ _0490_ _0493_ _0459_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout84_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3297_ _0424_ _0426_ _0427_ _0346_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4643__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4159__A1 Control_Unit.cont\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput34 net34 X[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput23 net23 X[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput45 net45 X[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4331__A1 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3437__A3 Control_Unit.T\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2948__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3070__A1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4570__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3220_ Control_Unit.T\[14\] _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3151_ _0289_ _0293_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3082_ _2112_ _0225_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2636__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3984_ _1050_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2935_ _2260_ _2261_ _2262_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2866_ _2176_ _1877_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4605_ _1976_ _1978_ _1979_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2797_ _2123_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4536_ _1558_ _1562_ _1379_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4467_ _1478_ _1474_ _1486_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3418_ Control_Unit.Q\[0\] Control_Unit.T\[0\] _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4398_ _2010_ _1403_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3349_ _0462_ _0463_ _0476_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2627__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2943__B _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3052__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3774__B _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2866__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2618__B2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3291__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2720_ _2040_ _1755_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2651_ _1976_ _1977_ _1978_ _1979_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2582_ _1792_ _1910_ _1827_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3346__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4321_ Control_Unit.Mc _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4693__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ _1303_ _1304_ _0841_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout109 net117 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3203_ _0339_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4183_ _1239_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2747__C _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3134_ Control_Unit.T\[0\] _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3065_ _0204_ _0205_ _0207_ _0210_ Control_Unit.futuro\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_27_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3034__A1 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3967_ _1018_ _1023_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_17_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2918_ _1913_ _2244_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3898_ _1798_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2849_ _2177_ _1966_ _1733_ _2173_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4534__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4519_ _1728_ _1534_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3025__B2 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3523__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3264__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3821_ _0832_ _0886_ _0834_ _0900_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3567__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3752_ _0821_ _0825_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2703_ _1727_ _1876_ _2028_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3683_ _0767_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2634_ _1888_ _1892_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2565_ _1866_ _1893_ _1862_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4304_ _0338_ Control_Unit.Mc _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2496_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4235_ _1287_ _1289_ _1290_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4166_ _1201_ _1207_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3117_ _0252_ _0256_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4097_ _0320_ _1148_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3048_ _1888_ _2317_ _0193_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3255__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3558__A2 _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3730__A2 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3494__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3246__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4174__I Control_Unit.Q\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3797__A2 Control_Unit.C\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout91 net94 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout80 net81 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2350_ Control_Unit.presente\[2\] _1677_ _1683_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4020_ _1075_ _1076_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3485__A1 _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2996__B1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3804_ net38 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4784_ _0108_ net67 Control_Unit.C\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3735_ net34 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3666_ _0749_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3597_ Control_Unit.T\[12\] _2019_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2617_ net13 _1945_ _1912_ _1909_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2548_ _1876_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3712__A2 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4218_ _0788_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2479_ _1807_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3476__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4149_ _1197_ _1198_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3228__A1 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3400__A1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2754__A3 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4754__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3219__A1 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4416__B1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3520_ _0617_ _0620_ _0539_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3451_ _2016_ Control_Unit.T\[2\] _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2402_ _1727_ _1730_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3382_ _2153_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4003_ _1029_ _1032_ _1048_ _1051_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4186__A2 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ _0091_ net90 Control_Unit.Q\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3718_ _0801_ _0803_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4698_ _0033_ net54 Control_Unit.cont\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4777__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2997__I _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3649_ _0734_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2415__A2 _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2951_ _2277_ _2278_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4168__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2882_ _1749_ _1895_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4621_ _1630_ _1631_ _1632_ _1634_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4552_ _0384_ _1988_ _1993_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4483_ _1420_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3503_ _0578_ _0590_ _0591_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3434_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3365_ _0468_ _0469_ _0491_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3296_ _0433_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout77_I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4159__A2 Control_Unit.Q\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4819_ _0143_ net61 Control_Unit.T\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 net24 X[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 X[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput46 net46 X[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4331__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3842__A1 Control_Unit.Q\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4398__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3070__A2 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2430__I _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3150_ _0289_ _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3081_ Control_Unit.T\[9\] _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2636__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2605__I _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3983_ _1029_ _1032_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3061__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2934_ _2144_ _2252_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2865_ _2191_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4604_ _1996_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4535_ _1559_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2796_ _2081_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2572__A1 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4466_ _1489_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3417_ _2014_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4815__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _1426_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3348_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3279_ _0415_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4001__A1 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2563__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3081__I Control_Unit.T\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2618__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2425__I _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3043__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2650_ Control_Unit.C\[26\] _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2554__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3256__I _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2581_ _1785_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4320_ _2014_ _2153_ _1359_ _1361_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4251_ _0936_ _1302_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3202_ _0327_ _0337_ _0341_ _0344_ _0345_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA_input1_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4182_ _1734_ _1219_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4059__A1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3133_ _0276_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3064_ _2025_ _0209_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_27_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3282__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4231__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3966_ _1016_ _1035_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2917_ _2241_ _2243_ _2242_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2793__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3897_ _1820_ _0967_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_13_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2848_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2779_ _2105_ _2085_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4518_ _1880_ Control_Unit.C\[15\] _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4449_ _2036_ _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4298__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3273__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2784__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2536__A1 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3804__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4289__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4461__A1 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3820_ _0893_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3751_ _0807_ _0811_ _0818_ _0826_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_14_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2702_ _1880_ _2030_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3567__A3 Control_Unit.Q\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3682_ _0768_ _0769_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2633_ net7 _1961_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2564_ _1851_ _1855_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_12_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4303_ _1344_ _1346_ _1347_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2495_ Control_Unit.cont\[4\] _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4234_ _0797_ _1274_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _1222_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3116_ _0259_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4096_ _1142_ _1147_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3047_ _1700_ _0189_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2766__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3558__A3 Control_Unit.Q\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3949_ _1796_ _0584_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_17_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4443__A1 _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout92 net93 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_35_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2757__A1 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout81 net88 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout70 net75 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_14_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3485__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3237__A2 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4434__A1 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2996__B2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2996__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3803_ _0872_ _0874_ _0882_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2748__A1 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ _0107_ net87 Control_Unit.Q\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3734_ _0725_ _0806_ _0727_ _0819_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3665_ _0744_ _0747_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2616_ _1942_ _1944_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3596_ _0361_ Control_Unit.C\[13\] Control_Unit.Q\[13\] _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2547_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2478_ _1802_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2920__A1 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4217_ _0950_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3476__A2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4148_ _0383_ _1208_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_44_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4079_ _1123_ _1124_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2523__I _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2911__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4416__A1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4134__B _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3450_ _0540_ _0553_ _0554_ _0555_ _0519_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_6_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3155__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2401_ _1728_ _1729_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3381_ _0503_ _0504_ _0505_ _0502_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2902__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4002_ _1067_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4095__I Control_Unit.Q\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4407__A1 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2608__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4766_ _0090_ net73 Control_Unit.Q\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3717_ _0801_ _0803_ _0776_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4697_ _0032_ net54 Control_Unit.cont\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3648_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3579_ net22 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3385__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3137__A1 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4637__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2428__I Control_Unit.cont\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2950_ _2240_ _2246_ _2267_ _2271_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_16_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2881_ _2208_ _1750_ _1865_ _1754_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _1379_ _1633_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4551_ _1569_ _1572_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4482_ _1505_ _1501_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3502_ _0600_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3433_ _0521_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3364_ Control_Unit.T\[28\] _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3295_ _0429_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3851__A2 Control_Unit.C\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4818_ _0142_ net61 Control_Unit.T\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4749_ _0073_ net97 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput25 net25 X[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput36 net36 X[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput47 net47 X[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3070__A3 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3080_ _1746_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4767__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3982_ _1025_ _1028_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2933_ _1927_ _1919_ _1921_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2864_ _2188_ _2189_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3349__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4603_ _1618_ _1616_ _1619_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2795_ _2080_ _2071_ _2079_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4534_ _0388_ _1542_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4465_ _1489_ _1487_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3416_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4396_ _1427_ _1432_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3347_ Control_Unit.T\[26\] _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3278_ _0416_ _0396_ _0410_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3824__A2 Control_Unit.C\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2531__I _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3760__A1 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3028__B1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2580_ net12 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3751__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4250_ _1297_ _1033_ _1300_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4181_ _1735_ _1234_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3201_ Control_Unit.T\[12\] _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3503__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3132_ _0274_ _0275_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4059__A2 Control_Unit.Q\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3063_ _1704_ _1972_ _0208_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4231__A2 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3965_ _1029_ _1032_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2916_ _2241_ _2242_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3896_ _1796_ _0964_ _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_17_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2847_ _2027_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2778_ _2106_ _2087_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4517_ _2026_ Control_Unit.C\[16\] _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4448_ _1123_ Control_Unit.C\[11\] _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4278__I Control_Unit.Q\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4379_ _1413_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3258__B1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4222__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2784__A2 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2536__A2 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2436__I _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3750_ _0523_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2701_ _1856_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3972__A1 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3681_ _0430_ _1992_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _1740_ _1884_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2563_ _1890_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4302_ _0976_ _1343_ Control_Unit.Q\[31\] _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4233_ _0947_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ _1799_ _1806_ _1818_ _1822_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4164_ _2027_ _1206_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4095_ Control_Unit.Q\[13\] _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3115_ _0251_ _0257_ _0258_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3046_ _2324_ _0188_ _0190_ _0191_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_fanout52_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4204__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3948_ _2255_ _1007_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3879_ _1811_ Control_Unit.Q\[1\] _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4140__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4443__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout60 net76 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout71 net74 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout82 net84 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout93 net94 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4198__A1 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3802_ _0872_ _0874_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4782_ _0106_ net86 Control_Unit.Q\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3733_ _0812_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3945__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3664_ _0728_ _0733_ _0740_ _0748_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2615_ _1833_ _1943_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3595_ net23 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2546_ _1743_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2920__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2477_ _1805_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4216_ _1266_ _1270_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4122__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4147_ _1201_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4078_ _2208_ _1140_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3029_ _1927_ _1688_ _0174_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3635__I _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4361__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2911__A2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4664__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3303__C _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3219__A3 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2427__A1 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4416__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _1710_ _1725_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4352__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _0503_ _0459_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4104__A1 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ _1768_ _1046_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2418__A1 Control_Unit.cont\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4407__A2 Control_Unit.C\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _0089_ net73 Control_Unit.Q\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3918__A1 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3716_ _0786_ _0792_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4696_ _0031_ net52 Control_Unit.cont\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3647_ _0735_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3578_ _0662_ _0663_ _0674_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4343__A1 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2529_ Control_Unit.cont\[8\] Control_Unit.cont\[9\] _1721_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4673__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2409__A1 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3082__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3385__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3137__A2 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4334__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3073__A1 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2880_ _2047_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4573__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4550_ _1993_ _1570_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _1506_ _1511_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4696__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3501_ _0584_ _0601_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3432_ _0529_ _0530_ _0524_ _0538_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3128__A2 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3363_ _0476_ _0487_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2887__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3294_ _0430_ _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2811__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0141_ net67 Control_Unit.T\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4748_ _0072_ net101 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4679_ _0014_ net110 Control_Unit.T\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput37 net37 X[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput26 net26 X[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput48 net48 X[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4619__A2 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2802__B2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3309__B _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3095__I _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4307__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2439__I _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3294__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3981_ _1048_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3597__A2 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2932_ _1916_ _1934_ _1809_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_16_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2863_ _2045_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3349__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2794_ net14 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4602_ _1978_ _1379_ _1615_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4533_ _1546_ _1547_ _1545_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4464_ _1490_ _1495_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3415_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4395_ _1429_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ Control_Unit.T\[24\] _0474_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3277_ _0387_ _0391_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3037__B2 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3588__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2812__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4474__I _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3028__A1 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3028__B2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4180_ Control_Unit.cont\[15\] _1238_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3200_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3131_ _2255_ _0264_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3267__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3062_ _1683_ _1678_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4384__I _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3019__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3964_ _1029_ _1032_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3895_ Control_Unit.cont\[1\] _1770_ Control_Unit.Q\[3\] _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2915_ _1943_ _1834_ _1788_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2846_ _1967_ _2173_ _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4519__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2777_ _2052_ _2105_ _2049_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4516_ _1543_ _1539_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4447_ _1468_ _1470_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4378_ _1784_ _1414_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3329_ _0457_ Control_Unit.T\[23\] _0451_ _0452_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_24_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3258__A1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3249__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2700_ _2028_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3972__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3680_ Control_Unit.T\[18\] _1992_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2631_ _1888_ _1892_ _1955_ _1958_ _1959_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2562_ _1744_ _1872_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3283__I Control_Unit.Rc vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4301_ Control_Unit.Q\[31\] _0936_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ _1286_ _1279_ _1282_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2493_ _1821_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ _1203_ _1205_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4094_ _0939_ _1153_ _1156_ _1112_ _1157_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3114_ _0250_ _0247_ _0249_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3045_ _1695_ _2321_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3947_ _1004_ _1006_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3458__I _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2362__I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3878_ _0944_ _0949_ _0952_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2829_ _2132_ _2157_ _2122_ _2126_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3715__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3403__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout72 net73 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout61 net66 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout83 net84 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_31_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2693__A2 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3642__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4198__A2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3801_ _0880_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _0105_ net83 Control_Unit.Q\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3732_ _0813_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3663_ net28 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2614_ _1843_ _1841_ _1786_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3594_ _0623_ _0675_ _0625_ _0689_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2545_ _1873_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2476_ _1802_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4215_ _1264_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4146_ _1710_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ _1122_ _1125_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3028_ _2274_ _2141_ _1687_ _1920_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2372__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2911__A3 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3624__A1 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2427__A2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4352__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4000_ _1040_ _1045_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3615__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4764_ _0088_ net72 Control_Unit.Q\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3715_ _0787_ _0791_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4695_ _0030_ net52 Control_Unit.cont\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3646_ _0714_ _0736_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2354__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4818__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__A2 Control_Unit.C\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3577_ _0668_ _0671_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2528_ _1716_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2459_ _1784_ _1787_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2657__A2 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4129_ _1882_ _1169_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__A2 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2550__I _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2593__A1 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4334__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3137__A3 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3073__A2 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3500_ _0254_ _2007_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4480_ _1508_ _1510_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3431_ _0534_ _0535_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4325__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3362_ _0338_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3293_ _0424_ _0426_ _0346_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3836__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2635__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4816_ _0140_ net68 Control_Unit.T\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4013__A1 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4747_ _0071_ net102 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4678_ _0013_ net110 Control_Unit.T\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3629_ _0706_ _0720_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput38 net38 X[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput27 net27 X[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput49 net49 X[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4790__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2545__I _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2802__A2 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4307__A2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4491__A1 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3046__A2 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3980_ _1036_ _1037_ _1047_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_44_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2931_ _2254_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2862_ _2188_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4601_ _1978_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2793_ net15 _2120_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_15_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ _1728_ _1987_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4463_ _1492_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3414_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _1765_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3345_ _0475_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout75_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3276_ _0414_ _0405_ _0408_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3809__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4234__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2796__A1 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2720__A1 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4686__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3130_ _0271_ _0273_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3061_ _0206_ _2185_ _2186_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3963_ _0938_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2914_ _1840_ _1845_ _1793_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3894_ _1802_ _0965_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2845_ _1727_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4515_ _1531_ _1536_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2776_ _2058_ _2084_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4446_ _1478_ _1474_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2950__A1 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4377_ _2073_ _2006_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2702__A1 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3328_ _0456_ _0458_ _0460_ _0455_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3259_ Control_Unit.T\[16\] _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4207__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3430__A2 Control_Unit.Q\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2941__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3603__B _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3249__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2630_ net5 _1957_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2561_ _1873_ _1889_ _1875_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2932__A1 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2492_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4300_ _1342_ _1344_ _1345_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4231_ _1279_ _1282_ _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4162_ _1706_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4093_ Control_Unit.Q\[12\] _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3113_ _0252_ _0256_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3044_ net5 _0189_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3946_ _0599_ _0951_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2620__B1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3877_ _0544_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2828_ _2137_ _2140_ _2156_ _2136_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2759_ _2058_ _2084_ _2085_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4429_ _1438_ _1440_ _1450_ _1460_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_8_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2553__I _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout73 net74 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_35_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout62 net66 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout95 net118 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout84 net86 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3333__B _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2693__A3 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4780_ _0104_ net83 Control_Unit.Q\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3800_ _0876_ _0879_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ _0814_ _0815_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3662_ _0662_ _0742_ _0752_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3593_ _0682_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2613_ _1823_ _1829_ _1836_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2544_ _1738_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2475_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4214_ _1245_ _1259_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4339__B _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4145_ _1203_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2638__I _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3330__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ _1122_ _1125_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_36_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3027_ _2274_ _2141_ _1937_ _1920_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3397__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3929_ _0985_ _0987_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3149__A1 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2372__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4649__A1 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3321__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3388__A1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4763_ _0087_ net72 Control_Unit.Q\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3714_ _0796_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4694_ _0029_ net52 Control_Unit.cont\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3645_ _0385_ _2020_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4343__A3 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3576_ _0668_ _0671_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2527_ _1742_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2458_ _1786_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2368__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2389_ Control_Unit.cont\[7\] _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2657__A3 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3854__A2 Control_Unit.C\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4128_ _1163_ _1168_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input18_I start vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4059_ _1714_ Control_Unit.Q\[11\] _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3199__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2593__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2741__I _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3430_ Control_Unit.C\[1\] Control_Unit.Q\[1\] _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3361_ _0442_ _0488_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3533__A1 Control_Unit.T\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3292_ Control_Unit.T\[18\] _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3049__B1 _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4815_ _0139_ net87 Control_Unit.C\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ _0070_ net103 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3772__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4677_ _0012_ net92 Control_Unit.T\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3628_ _0707_ _0710_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput39 net39 X[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput28 net28 X[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3559_ Control_Unit.T\[9\] Control_Unit.C\[9\] _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4619__A4 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3515__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3392__I _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4808__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2930_ _2133_ _2257_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2861_ _1740_ _1875_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4600_ _1616_ _1617_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2792_ net16 _2114_ _2120_ _1689_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4531_ _1550_ _1555_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4462_ _0224_ _2003_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3506__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3413_ _0520_ Control_Unit.Mx _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4393_ _1831_ Control_Unit.C\[7\] _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3344_ _0473_ _0466_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3275_ _0404_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4482__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout68_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4234__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3993__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2381__I _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4729_ _0053_ net78 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2720__A2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__B _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3276__A3 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output49_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4161__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3060_ _1702_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3962_ _1030_ _1012_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2913_ _1840_ _1845_ _1792_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3893_ _1803_ Control_Unit.Q\[2\] _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2844_ _1874_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3727__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4514_ _1989_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2775_ _2103_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4445_ _1477_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2950__A2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4376_ _2073_ Control_Unit.C\[5\] _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2702__A2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3327_ _0456_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3258_ _0380_ _0393_ _0396_ _0397_ _0398_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__3258__A3 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2376__I _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3189_ _0312_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2769__A2 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4391__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2941__A2 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4143__A1 Control_Unit.cont\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout118_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2560_ _1735_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4382__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2932__A2 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2491_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4134__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4230_ _1283_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4161_ _1218_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4092_ _1138_ _1154_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3112_ _0245_ _0253_ _0255_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3043_ _2220_ _2302_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4625__B _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3948__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3945_ _0996_ _1013_ _1015_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2620__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3876_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2827_ _1703_ _2139_ _2142_ _1687_ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2758_ _2086_ _2048_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4676__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4125__A1 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2689_ Control_Unit.C\[13\] _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4428_ _1364_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__I _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4359_ _2008_ _0971_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout74 net75 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout63 net65 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net54 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout85 net86 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout96 net100 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2914__A2 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2744__I _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ _0445_ _1981_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2602__A1 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4699__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3661_ _0748_ _0750_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3575__I _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3592_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2612_ _1909_ _1912_ _1924_ net11 _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2543_ _1745_ _1871_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4107__A1 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2474_ _1770_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4658__A2 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2669__A1 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4144_ _1712_ _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3330__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4075_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3026_ _1931_ _1930_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2654__I Control_Unit.C\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3397__A2 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4594__A1 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3928_ _0979_ _0997_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3859_ _0540_ _0933_ _0934_ _0935_ _0582_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4346__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2372__A3 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4649__A2 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2832__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2899__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3560__A2 Control_Unit.C\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4762_ _0086_ net71 Control_Unit.Q\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3379__A2 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _0797_ _0798_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4693_ _0028_ net52 Control_Unit.cont\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3644_ _0385_ _2020_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3575_ _0522_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2526_ _1853_ _1854_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_fanout98_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2649__I Control_Unit.C\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2457_ _1785_ _1772_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2388_ Control_Unit.cont\[6\] _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__2657__A4 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ _0388_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4058_ _1715_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3009_ _2267_ _2271_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4567__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4319__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3943__I _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3542__A2 Control_Unit.C\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2559__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2750__B1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2805__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3339__B _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout100_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4737__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3360_ _0462_ _0463_ _0476_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2469__I _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3291_ _0422_ _0428_ _0342_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4814_ _0138_ net84 Control_Unit.C\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _0069_ net103 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4676_ _0011_ net92 Control_Unit.T\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3772__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3627_ _0711_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3558_ Control_Unit.T\[10\] _2004_ Control_Unit.Q\[10\] _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xoutput29 net29 X[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2379__I _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2509_ _1776_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3489_ _0590_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3288__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3460__A1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3451__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2860_ _1881_ _1876_ _1890_ _2030_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2791_ _2117_ _2119_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_15_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4530_ _1988_ _1354_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4461_ _2036_ _1481_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3506__A2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3412_ Control_Unit.Rx _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4392_ _1910_ _1405_ _1428_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ Control_Unit.T\[25\] _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3274_ Control_Unit.T\[17\] _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__4628__B _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2927__I _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3690__A1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3442__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2662__I _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2989_ _2303_ _2316_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4728_ _0052_ net79 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ _0306_ _0259_ _0330_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3681__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4704__D _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3672__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3961_ _0999_ _1009_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2912_ _1793_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2482__I _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3892_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2843_ _2094_ _2170_ _2171_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2774_ net7 _2099_ _2102_ net6 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3727__A2 Control_Unit.C\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4513_ _1538_ _1540_ _1541_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4202__I _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4444_ _1466_ _1471_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4375_ _1838_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3326_ _0375_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout80_I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3257_ _0385_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3188_ _0329_ _0331_ _0309_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4022__I _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2932__A3 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2490_ _1769_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3861__I _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4160_ _1709_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2477__I _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3111_ _0254_ _1826_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _1152_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3042_ _1696_ _2323_ _0153_ _0186_ _0187_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_23_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3944_ _0584_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3101__I _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3875_ _0945_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2826_ _2154_ _2146_ _2147_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2620__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2757_ _2030_ _1750_ _2038_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2688_ _2013_ _2014_ _2015_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4427_ _2000_ _1407_ _1436_ _1461_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3884__A1 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4358_ _1831_ _1820_ _2006_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3309_ _0422_ _0439_ _0343_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4289_ _0490_ _1336_ _0950_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4061__A1 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout53 net54 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout75 net76 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout97 net100 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout86 net87 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2375__A1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4770__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3630__B _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4052__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2602__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3660_ _0748_ _0750_ _0672_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3591_ _0683_ _0686_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2611_ _1936_ _1938_ _1939_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2542_ _1867_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4212_ Control_Unit.Q\[19\] _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2473_ _1801_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3866__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2669__A2 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4143_ Control_Unit.cont\[12\] Control_Unit.Q\[15\] _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4074_ _1128_ _1131_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4636__B _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3025_ _1692_ _0165_ _0170_ _1693_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4043__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3927_ _0982_ _0988_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3858_ net43 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3789_ _0832_ _0859_ _0834_ _0870_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2809_ _1913_ _1806_ _2074_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2372__A4 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2845__I _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4034__A1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4712__D _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__A2 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3388__A3 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2580__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2520__A1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ _0085_ net56 Control_Unit.Q\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3712_ Control_Unit.T\[20\] _1983_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4692_ _0027_ net99 Control_Unit.T\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3643_ _0399_ Control_Unit.C\[16\] Control_Unit.Q\[16\] _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4328__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3574_ _0655_ _0669_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2525_ _1759_ _1781_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2456_ _1773_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _1182_ _1187_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2387_ Control_Unit.cont\[10\] _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2511__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4366__B _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4264__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _1718_ _1113_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3008_ _2267_ _2271_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4567__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__A2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3445__B _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2750__A1 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4689__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4276__B _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3290_ _0424_ _0426_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4549__A2 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4813_ _0137_ net85 Control_Unit.C\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4744_ _0068_ net102 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4675_ _0010_ net90 Control_Unit.T\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3626_ _0715_ _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 net19 X[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3557_ _0650_ _0654_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2508_ _1833_ _1836_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3488_ _0585_ _0589_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4485__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3288__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2439_ _1767_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109_ _1159_ _1160_ _1170_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_5_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2799__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3460__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4115__I Control_Unit.Q\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2971__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2723__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4476__A1 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4228__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3451__A2 Control_Unit.T\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4704__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2790_ _2118_ _2082_ _2065_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__I _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _2041_ _1491_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2962__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3411_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4391_ _1839_ _1412_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2714__A1 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3342_ _0377_ _0465_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3273_ _0399_ _0363_ _0411_ _0412_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_6_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4219__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3442__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2988_ _2309_ _2315_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4727_ _0051_ net78 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4658_ _0231_ _1644_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3609_ _0691_ _0694_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2705__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _1356_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3681__A2 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2944__A1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4449__A1 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ _0999_ _1009_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2911_ _2063_ _1904_ _2238_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_16_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3891_ _1810_ Control_Unit.Q\[2\] _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2842_ _2029_ _2096_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2773_ _2091_ _2101_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4512_ _2020_ _1403_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _2004_ _1462_ _1474_ _1476_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4374_ _1824_ Control_Unit.C\[6\] _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3325_ _0445_ _0457_ _0378_ _0439_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3360__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3256_ _0343_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3112__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3187_ _0259_ _0330_ _0306_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__D _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3179__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2848__I _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3351__A1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3103__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3654__A2 Control_Unit.C\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4715__D _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3590__A1 Control_Unit.Q\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3342__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3110_ Control_Unit.T\[5\] _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _1135_ _1110_ _1132_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3645__A2 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3041_ _2325_ _2331_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2493__I _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3943_ _0950_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3874_ _0947_ _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2825_ _2153_ net2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4213__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2908__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2756_ _2049_ _2052_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2687_ Control_Unit.C\[2\] _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4426_ _1454_ _1460_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2668__I Control_Unit.C\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3333__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4357_ _1388_ _1390_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3308_ _0442_ _0439_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4288_ _1332_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3239_ _0346_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout65 net66 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout54 net55 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout76 net119 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout87 net88 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2375__A2 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3590_ Control_Unit.Q\[11\] _0684_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2610_ net11 _1924_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2541_ _1869_ _1862_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3872__I _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2472_ _1800_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4211_ _1707_ _0768_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3315__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2669__A3 Control_Unit.C\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4142_ _1713_ _1177_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4073_ _1114_ _1115_ _1134_ _1137_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3024_ _2276_ _0169_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4043__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3926_ _0982_ _0988_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3857_ _0926_ _0932_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3788_ _0864_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2808_ _1909_ _2135_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2357__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2739_ _1787_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3554__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3306__B2 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3306__A1 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4409_ _1832_ Control_Unit.C\[7\] _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3609__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2348__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3545__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _0084_ net56 Control_Unit.Q\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3711_ Control_Unit.T\[20\] Control_Unit.C\[20\] _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4691_ _0026_ net96 Control_Unit.T\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3642_ _0728_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3536__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3573_ _0656_ _0659_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2524_ _1852_ _1753_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2455_ _1783_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2386_ Control_Unit.cont\[9\] _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3839__A2 Control_Unit.C\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4125_ _1735_ _1184_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2946__I _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4056_ _1752_ _1101_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3007_ _2325_ _2331_ _2334_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3777__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4813__D _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2681__I Control_Unit.C\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3909_ _0965_ _0968_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3527__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2591__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3687__I _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4191__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4783__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4812_ _0136_ net84 Control_Unit.C\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4743_ _0067_ net102 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4674_ _0009_ net89 Control_Unit.T\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3625_ Control_Unit.Q\[14\] _0716_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4182__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3556_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2507_ _1826_ _1835_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3487_ _0585_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2438_ _1766_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2369_ net16 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4808__D _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4108_ _1159_ _1160_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4039_ _1079_ _1085_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input16_I n[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4131__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2723__A2 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__A1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4306__I _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3366__B _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2962__A2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4164__A1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3410_ Control_Unit.Mx _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4390_ _1413_ _1416_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2714__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3341_ _0472_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3272_ _0402_ _0410_ _0378_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input8_I n[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3675__B1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2496__I _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3978__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2987_ _2308_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2402__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4726_ _0050_ net78 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4679__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4657_ _0341_ _1660_ _1661_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4155__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3608_ _0691_ _0694_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2705__A2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4588_ _1607_ _1606_ _1604_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3539_ _0623_ _0624_ _0625_ _0638_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4630__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4570__B _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2944__A2 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4146__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2632__A1 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2910_ _1845_ _1792_ _1849_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3890_ _0960_ _0962_ _0963_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2841_ _2029_ _2096_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2772_ _2100_ _2090_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4511_ _1422_ _1539_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4137__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4442_ _1422_ _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2699__A1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4373_ _1397_ _1400_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3324_ Control_Unit.T\[22\] _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3360__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3255_ _0381_ _0394_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout66_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3186_ _0261_ _0269_ _0301_ _0304_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2871__A1 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2623__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2623__B2 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3179__A2 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__A1 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4709_ _0152_ _4709_/E _4709_/RN Control_Unit.Rc vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__4128__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3103__A2 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output47_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4119__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2696__A4 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3040_ _0163_ _0178_ _0179_ _0185_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2853__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3942_ _0999_ _1009_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3873_ _1813_ _0531_ _0943_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2824_ _1928_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4358__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2755_ _2060_ _2061_ _2062_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2686_ Control_Unit.C\[3\] _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4425_ _1447_ _1459_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4717__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4356_ _1382_ _1387_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3333__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3307_ _0376_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4287_ _1334_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3238_ _0362_ _0363_ _0373_ _0379_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3097__A1 _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3169_ _0236_ _0311_ _0312_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout55 net60 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout99 net100 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout66 net70 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout88 net95 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout77 net80 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3088__A1 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4052__A3 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__I _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout116_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2540_ _1868_ _1859_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2471_ Control_Unit.cont\[1\] _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4210_ _1256_ _1257_ _1255_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4512__A1 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4141_ _1736_ _1185_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4072_ _1135_ _1110_ _1132_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3079__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3023_ _2275_ _0168_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__B1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4579__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3925_ _0939_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _0926_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3787_ _0839_ _0865_ _0868_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2807_ _1692_ _2130_ _2135_ _1909_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2738_ _1717_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3554__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2679__I Control_Unit.C\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4503__A1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4408_ _2059_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2669_ _1995_ _1996_ Control_Unit.C\[31\] _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4339_ _1371_ _1378_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2817__A1 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3490__A1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3545__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3710_ Control_Unit.Q\[20\] _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _0025_ net85 Control_Unit.T\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3784__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3641_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3572_ _0660_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2523_ _1715_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2454_ _1774_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2385_ Control_Unit.cont\[8\] _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4124_ _1711_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 clk net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2448__B _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4055_ _1852_ _1118_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3006_ _1698_ _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3472__A1 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3908_ _0965_ _0968_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3839_ _0497_ Control_Unit.C\[30\] Control_Unit.Q\[30\] _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3527__A2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3463__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4191__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3208__I _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3454__A1 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2782__I _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ _0135_ net99 Control_Unit.C\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4742_ _0066_ net101 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4673_ _0008_ net89 Control_Unit.T\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3624_ _0366_ _2021_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3555_ _0645_ _0651_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout96_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3486_ _0586_ _0587_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2506_ _1834_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2437_ _1765_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2368_ net17 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4107_ _1889_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4038_ _0215_ _1098_ _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2692__I Control_Unit.C\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4173__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3739__A2 Control_Unit.C\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4322__I _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3911__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3340_ _0466_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3271_ _0402_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3675__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3675__B2 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3427__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2986_ _2207_ _2310_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_33_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4725_ _0049_ net78 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2461__B _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4656_ _0240_ _1642_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4155__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3607_ _0676_ _0681_ _0688_ _0695_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4587_ _1603_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3538_ _0631_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2687__I Control_Unit.C\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3469_ _0540_ _0567_ _0572_ _0573_ _0519_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3467__B _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4082__A1 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3221__I _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2632__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2840_ net8 _2097_ _2104_ _2168_ _2099_ _1964_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2396__A1 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2771_ _2039_ _2043_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _1530_ _1527_ _1537_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4441_ _1463_ _1465_ _1473_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4372_ _1408_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3323_ Control_Unit.T\[23\] _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3254_ _0392_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3185_ _0244_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout59_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2969_ _2289_ _2292_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4708_ _0043_ net90 Control_Unit.cont\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4796__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _0270_ _1644_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4064__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2880__I _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3660__B _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4055__A1 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4047__I Control_Unit.Q\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3941_ _1010_ _0994_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_17_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3872_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2823_ _2121_ _2122_ _2151_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4358__A2 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2754_ _2066_ _2069_ _2081_ _2082_ _2056_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_9_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2685_ Control_Unit.C\[0\] _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4424_ _1456_ _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3869__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4355_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3306_ _0344_ _0440_ _0441_ _0438_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4286_ _1333_ _1316_ _1325_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3237_ _0374_ _0360_ _0371_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3097__A2 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3168_ _0223_ _0228_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3099_ _0238_ _0241_ _0242_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2914__B _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout56 net60 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout89 net90 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout67 net69 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout78 net80 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3745__B _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2780__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4811__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3260__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout109_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2470_ _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ _1879_ _1199_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3079__A2 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _0946_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4276__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3022_ _0167_ _2262_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3924_ _0586_ _0937_ _0940_ _0995_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3251__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3539__B1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3855_ _0930_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3786_ _0850_ _0853_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2806_ _2068_ _2133_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_30_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2737_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2668_ Control_Unit.C\[30\] _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4407_ _1838_ Control_Unit.C\[8\] _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2599_ _1921_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2514__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _1348_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4269_ _1306_ _1317_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2817__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4019__A1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2538__C _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _0721_ _0730_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ _0664_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2522_ _1756_ _1764_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2453_ _1781_ _1778_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2384_ Control_Unit.cont\[11\] _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_25_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4123_ Control_Unit.cont\[11\] Control_Unit.Q\[14\] _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4054_ _1100_ _1102_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput2 n[0] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_3005_ _2329_ _2332_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_37_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3472__A2 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4421__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3907_ _1910_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3838_ _0907_ _0914_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3769_ Control_Unit.T\[24\] _1977_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3463__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4479__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3454__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4810_ _0134_ net98 Control_Unit.C\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _0065_ net101 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4672_ _0316_ _0347_ _1671_ _0397_ _1672_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3623_ Control_Unit.T\[14\] _2021_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3554_ _0640_ _0643_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3390__A1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3485_ _0262_ _2009_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2505_ _1827_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2436_ _1760_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout89_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2367_ net3 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4106_ _1163_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4037_ _1746_ _1100_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_25_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3445__A2 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2956__A1 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4330__B1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3684__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2947__A1 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3270_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2985_ _2199_ _2312_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4724_ _0048_ net77 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4655_ _1659_ _0304_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3606_ net24 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ _1977_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3537_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3468_ net44 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2419_ _1746_ _1747_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3399_ _0510_ _1863_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4579__B _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3354__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3106__A1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2617__B1 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2770_ _2093_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2396__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4440_ _1463_ _1465_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ _1394_ _1395_ _1401_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3322_ _0447_ _0344_ _0454_ _0455_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3253_ _0374_ _0360_ _0371_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3184_ _0229_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4073__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4243__I _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2968_ _2283_ _2287_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4707_ _0042_ net74 Control_Unit.cont\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2899_ _2118_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4638_ _1645_ _1647_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2698__I _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3336__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4399__B _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4569_ _1584_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4740__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3232__I _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ _0990_ _0992_ _0989_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ Control_Unit.Rc _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4358__A3 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2822_ _2132_ _2136_ _2150_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2753_ _2064_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2684_ Control_Unit.C\[1\] _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4423_ _2067_ _2001_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3869__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4354_ _1383_ _1386_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2541__A2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3305_ _0435_ _0434_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4285_ _0895_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3236_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3167_ _0244_ _0308_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3098_ _0239_ _0240_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4763__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout57 net58 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout79 net80 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4349__A3 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout68 net69 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3309__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4037__A2 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3987__I Control_Unit.Q\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3796__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4070_ _1116_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3079__A3 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4058__I _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3021_ _2260_ _2261_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3923_ _0989_ _0993_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3854_ _0503_ Control_Unit.C\[31\] Control_Unit.Q\[31\] _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3539__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2805_ _2074_ _2076_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3785_ _0855_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2736_ _1767_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2667_ Control_Unit.C\[28\] _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4406_ _1429_ _1431_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2598_ _1926_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4337_ _1367_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4268_ _1111_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3219_ _0347_ _0356_ _0360_ _0344_ _0361_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4267__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4199_ _1706_ _1238_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3950__A1 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3491__B _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3570_ Control_Unit.Q\[10\] _0665_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2521_ _1768_ _1780_ _1782_ _1847_ _1849_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_6_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2452_ _1762_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2383_ Control_Unit.cont\[13\] _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4122_ _0215_ _1158_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4053_ _1100_ _1102_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4249__A2 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3004_ _2273_ _2279_ _2288_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xinput3 n[10] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3906_ _0975_ _0977_ _0978_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3576__B _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2983__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4801__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3837_ _0902_ _0905_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4185__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3768_ Control_Unit.T\[24\] _1977_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2719_ _2047_ _1754_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3699_ _0438_ Control_Unit.C\[20\] Control_Unit.Q\[20\] _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4488__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__A1 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4660__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4100__A1 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2565__B _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2414__A1 Control_Unit.cont\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4740_ _0064_ net97 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4671_ _0213_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4167__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3622_ Control_Unit.T\[15\] Control_Unit.C\[15\] _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_30_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4071__I _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3914__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3553_ _0640_ _0643_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3484_ _0262_ _2009_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2504_ _1832_ _1791_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3390__A2 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2435_ _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3415__I _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4105_ _0351_ _1165_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2366_ net4 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ _1752_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2956__A2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4158__A1 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3905__A1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4330__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4094__B1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3060__I _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2947__A2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2984_ _2206_ _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4723_ _0047_ net67 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4654_ _0257_ _1657_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4585_ _1603_ _1357_ _1604_ _1605_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3605_ _0662_ _0690_ _0699_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3536_ _0632_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3467_ _0568_ _0569_ _0570_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4312__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2418_ Control_Unit.cont\[8\] _1722_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3398_ _0510_ _1864_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2874__A1 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2349_ Control_Unit.presente\[0\] _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4019_ _0224_ _1079_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_input14_I n[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4615__A2 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2626__B2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2626__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2933__B _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2929__A2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3051__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4551__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3106__A2 Control_Unit.T\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2617__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3042__A1 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3042__B2 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2396__A3 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4370_ _1394_ _1401_ _1390_ _1388_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3321_ _0447_ _0453_ _0442_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3896__A3 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3252_ _0382_ _0373_ _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3183_ _0221_ _0316_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_26_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input6_I n[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2967_ _2289_ _2292_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3033__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4706_ _0041_ net71 Control_Unit.cont\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2898_ _2222_ _2223_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4637_ _0281_ _0286_ _1646_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3336__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ _1588_ _1590_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_2_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _1349_ _1526_ _1527_ _1406_ _1528_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3519_ _0618_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4692__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3327__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2838__B2 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2838__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3870_ Control_Unit.Mq _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2821_ _2137_ _2140_ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_13_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2752_ _2071_ _2079_ _2080_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3318__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ _1759_ _1443_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2683_ _2007_ _2009_ _2010_ _2011_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4353_ _1350_ _1391_ _1392_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3304_ _0380_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4284_ Control_Unit.Q\[28\] _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3235_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3423__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3097_ _0239_ _0240_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4254__I Control_Unit.Q\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout58 net59 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3006__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3999_ _2060_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout69 net70 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4506__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output45_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3245__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3796__A2 Control_Unit.C\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2412__I _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3243__I _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3484__A1 _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3020_ _1692_ _0165_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3922_ _0970_ _0973_ _0974_ _0961_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_3853_ _0927_ _0928_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2804_ _1918_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3784_ _0850_ _0853_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2735_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2666_ Control_Unit.C\[29\] _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _1438_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3711__A2 Control_Unit.C\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2597_ _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4336_ _1373_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4267_ _1318_ _1316_ _1136_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4198_ _2026_ _0743_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3218_ Control_Unit.T\[13\] _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3475__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4672__B1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3149_ _1934_ _0291_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3227__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3778__A2 Control_Unit.C\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3702__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3466__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2407__I Control_Unit.cont\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3769__A2 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout114_I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2520_ _1848_ _1844_ _1842_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_10_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2451_ _1779_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2382_ Control_Unit.cont\[12\] _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4753__CLK net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4121_ _1868_ _1166_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4052_ _1088_ _1108_ _1096_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3457__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3003_ _2330_ _2293_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xinput4 n[11] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3209__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3905_ _0563_ _0951_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2432__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3836_ _0902_ _0905_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3767_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2718_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3932__A2 Control_Unit.Q\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3698_ _0780_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2649_ Control_Unit.C\[27\] _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4319_ _0525_ _0941_ _1359_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4645__B1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2936__B _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4176__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4776__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4598__B _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2414__A2 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ _0328_ _0334_ _0314_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3621_ Control_Unit.Q\[15\] _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3914__A2 Control_Unit.Q\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3552_ _0627_ _0630_ _0637_ _0644_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2503_ _1831_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3483_ Control_Unit.Q\[4\] _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2434_ _1758_ _1759_ _1762_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2365_ _1690_ _1691_ _1692_ _1693_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4104_ _1868_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ _1760_ Control_Unit.Q\[10\] _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3819_ _0894_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4799_ _0123_ net92 Control_Unit.C\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3905__A2 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4211__B _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2510__I _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2420__I _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4085__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3832__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2983_ _2207_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4722_ _0046_ net67 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4653_ _1657_ _0347_ _1658_ _0397_ _0598_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3604_ _0695_ _0697_ _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4584_ _1603_ _1601_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3535_ _0611_ _0633_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3466_ _0562_ _0564_ _0565_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2417_ Control_Unit.cont\[9\] _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3397_ _0510_ _1758_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2874__A2 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2348_ _1675_ _1682_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4018_ _2059_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2626__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2562__A1 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3106__A3 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3071__I _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3042__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3320_ _0447_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_4_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3690__B _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3251_ _0387_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3182_ _0321_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3805__B2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3805__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2966_ _2273_ _2279_ _2288_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4705_ _0040_ net58 Control_Unit.cont\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2897_ _2222_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2792__A1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2792__B2 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4636_ _0281_ _0286_ _0340_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4567_ _1588_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _2021_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3518_ _0604_ _0608_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3449_ net41 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3272__A2 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4221__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4460__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2820_ _1930_ _2143_ _2146_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2751_ _1779_ _1787_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2774__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2774__B2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2682_ Control_Unit.C\[6\] _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _1123_ _1455_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4352_ _2009_ _1354_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3303_ _0424_ _0426_ _0437_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_28_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4283_ _1331_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4279__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3234_ Control_Unit.Rc _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3165_ _0230_ _0234_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout57_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3096_ Control_Unit.T\[7\] _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A1 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout59 net60 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3998_ _1059_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2949_ _2240_ _2246_ _2276_ _1944_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4619_ _1627_ _1996_ _1997_ _1622_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_11_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2508__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3181__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3524__I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3484__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4433__A1 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4682__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3921_ _0990_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3852_ _0500_ Control_Unit.C\[30\] _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2803_ _2126_ _2131_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3783_ _0846_ _0854_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2734_ _1844_ _1842_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2665_ _1988_ _1989_ _1991_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2596_ _1807_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4404_ _1427_ _1425_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4335_ _1798_ _1374_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3434__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4266_ _1306_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4197_ _1706_ _1251_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3217_ _0357_ _0358_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3475__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3148_ _1926_ _0290_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3227__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3079_ _2050_ _0216_ _0222_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3778__A3 Control_Unit.Q\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2910__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2423__I _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2729__A1 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2450_ _1778_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout107_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2381_ _1709_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ _0319_ _1180_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4051_ _1104_ _1107_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_7_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3002_ _2296_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput5 n[12] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3904_ _0961_ _0974_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3429__I Control_Unit.T\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3835_ _0889_ _0892_ _0899_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3766_ Control_Unit.T\[25\] Control_Unit.C\[25\] Control_Unit.Q\[25\] _0849_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2717_ Control_Unit.cont\[10\] _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3393__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3697_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3145__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2648_ Control_Unit.C\[24\] _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2579_ _1846_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4318_ _1360_ _1809_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4249_ _1297_ _1112_ _1301_ _1302_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_28_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4636__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3620_ net25 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3551_ net20 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2502_ _1774_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3127__A1 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3482_ Control_Unit.T\[5\] _2006_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2433_ _1760_ _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2364_ net12 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4103_ _1716_ Control_Unit.Q\[13\] _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4034_ _1848_ _1074_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3818_ _0895_ _0896_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4798_ _0122_ net91 Control_Unit.C\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3366__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3749_ net35 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2629__B1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2644__A3 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3841__A2 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3109__A1 Control_Unit.T\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4609__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3688__B _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2982_ _2303_ _2308_ _2309_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4721_ _0045_ net77 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _0269_ _0301_ _0261_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3603_ _0695_ _0697_ _0672_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ _1588_ _1590_ _1599_ _1983_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3534_ _0240_ _2010_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3465_ _0561_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2416_ _1742_ _1743_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ _0512_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout87_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2347_ Control_Unit.presente\[2\] _1674_ _1681_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4017_ _1081_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4766__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3339__A1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2562__A2 _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3511__A1 Control_Unit.T\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3814__A2 Control_Unit.C\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3578__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2431__I Control_Unit.cont\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3250_ _0388_ _0389_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3181_ _0322_ _0323_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3502__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4789__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4093__I Control_Unit.Q\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4704_ _0039_ net71 Control_Unit.cont\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2965_ _2289_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2896_ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4635_ _0290_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _1543_ _1539_ _1589_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3741__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3517_ _0600_ _0603_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4497_ _1517_ _1515_ _1525_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3448_ _0548_ _0552_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4297__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ _0500_ _0378_ _0488_ _0498_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__B1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2750_ _2064_ _1835_ _2072_ _2078_ _2071_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2681_ Control_Unit.C\[7\] _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4420_ _1760_ Control_Unit.C\[9\] _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4351_ _1388_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3302_ Control_Unit.T\[20\] _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4282_ _0895_ _1329_ _1330_ _1317_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3233_ Control_Unit.Mt _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3164_ _0260_ _0305_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3095_ _1839_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4451__A2 _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2462__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4804__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ _0238_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2948_ _1829_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2879_ _2200_ _2205_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4618_ _1997_ _1403_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2517__A2 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4549_ _1565_ _1365_ _1573_ _1574_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_2_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3478__B1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3650__B1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3540__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4433__A2 Control_Unit.C\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4827__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3920_ _1822_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3851_ _0500_ Control_Unit.C\[30\] _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4197__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3782_ _0860_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2802_ _1691_ _2081_ _2124_ _2130_ net13 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2733_ _1755_ _1780_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2747__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3944__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2664_ _1992_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2595_ _1919_ _1923_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4403_ _1432_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4334_ _2016_ _1804_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4121__A1 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4265_ _0938_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4196_ _1247_ _1252_ _1253_ _1231_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3216_ _0355_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4672__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3147_ _1925_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3078_ _2208_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2986__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__A1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4360__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2910__A2 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output50_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4179__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2729__A2 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2380_ Control_Unit.cont\[14\] _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4103__A1 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ _1111_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3001_ _2326_ _2327_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput6 n[13] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3090__A1 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3903_ _0946_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3834_ _0906_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3917__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3765_ net36 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2716_ _1856_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3696_ _0773_ _0782_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3393__A2 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__A1 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2647_ Control_Unit.C\[25\] _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2578_ _1830_ _1837_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4317_ _2013_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ _1297_ _1300_ _1136_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4645__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4179_ _1734_ Control_Unit.Q\[17\] _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2408__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4581__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4333__A1 Control_Unit.C\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2895__A1 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3550_ _0582_ _0639_ _0648_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3375__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2501_ _1788_ _1794_ _1823_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3127__A2 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4324__A1 Control_Unit.C\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3481_ Control_Unit.Q\[5\] _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2432_ _1717_ _1719_ _1720_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2363_ net13 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4102_ _0224_ _1157_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4033_ _1765_ _1082_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4627__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3063__A1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4797_ _0121_ net89 Control_Unit.C\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3817_ _0484_ Control_Unit.C\[27\] _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4563__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3748_ _0528_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4695__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ Control_Unit.Q\[18\] _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3175__I _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2877__A1 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3903__I _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4618__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2629__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2629__B2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3054__A1 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4554__A1 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3109__A2 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2873__B _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2981_ _2306_ _2307_ _2304_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3045__A1 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4720_ _0044_ net77 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4651_ _0261_ _0269_ _0301_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4545__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3602_ _0682_ _0687_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4582_ _1984_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3533_ Control_Unit.T\[7\] _2010_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3464_ _0548_ _0552_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2415_ _1736_ _1742_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3395_ _0511_ _2118_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2346_ _1680_ _1681_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4016_ _1765_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3823__A3 Control_Unit.Q\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4222__C _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3633__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3511__A2 Control_Unit.C\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3814__A3 Control_Unit.Q\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3027__B2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3027__A1 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2712__I _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3180_ _0222_ _0213_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2561__I0 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3018__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2964_ _2082_ _2290_ _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_15_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3569__A2 Control_Unit.C\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4703_ _0038_ net57 Control_Unit.cont\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2895_ _1866_ _1753_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4518__A1 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4634_ _0375_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4565_ _1553_ _1562_ _1585_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3516_ _0613_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4496_ _1517_ _1515_ _1525_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3447_ _0548_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3378_ Control_Unit.T\[31\] _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I n[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4284__I Control_Unit.Q\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3009__A1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4221__A3 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3248__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2707__I _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2680_ _2008_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4350_ _1370_ _1366_ _1389_ _1377_ _1367_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3723__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3301_ _0430_ _0435_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4756__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4369__I _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4281_ _0895_ _1325_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3232_ _0364_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input4_I n[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3163_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3094_ _1718_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ _1061_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2947_ _2274_ _1920_ _1922_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2878_ _2200_ _2205_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4617_ _1627_ _1620_ _1623_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _1569_ _1572_ _1421_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3714__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4479_ _0215_ _1502_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3478__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4427__B1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2527__I _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3650__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3650__B2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3469__B2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3469__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3850_ Control_Unit.Q\[30\] _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4197__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3781_ Control_Unit.Q\[25\] _0861_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2801_ _2129_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2732_ _1778_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__3944__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2663_ Control_Unit.C\[18\] _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2594_ _1920_ _1806_ _1922_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4402_ _1408_ _1409_ _1437_ _1433_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4333_ Control_Unit.C\[2\] _1804_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4264_ _1311_ _1313_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3215_ _0221_ _0316_ _0326_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4195_ _1228_ _1248_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3146_ Control_Unit.T\[2\] _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3880__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout62_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2683__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3077_ _0220_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3632__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3178__I _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3979_ _1036_ _1037_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3699__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4360__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output43_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3871__A1 Control_Unit.Rc vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4103__A2 Control_Unit.Q\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3551__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3000_ _2282_ _2287_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput7 n[14] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3902_ _0961_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3833_ net42 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3764_ _0832_ _0833_ _0834_ _0847_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2715_ _2039_ _2043_ _2042_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3695_ _0767_ _0781_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2646_ net18 _1684_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4342__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2577_ _1689_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4316_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4247_ _1297_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4178_ _1222_ _1224_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3129_ _1822_ _0272_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2408__A2 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4292__I Control_Unit.Q\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3908__A2 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4581__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4817__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4333__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2895__A2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4097__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4572__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout112_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3480_ net46 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2500_ _1787_ _1826_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2431_ Control_Unit.cont\[7\] _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2886__A2 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2362_ net14 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4101_ _2047_ _1145_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4032_ _2111_ _1084_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3835__A1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4260__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3063__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2561__S _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _0120_ net73 Control_Unit.C\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3816_ _0484_ Control_Unit.C\[27\] _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3747_ _0765_ _0820_ _0831_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2360__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3678_ Control_Unit.T\[19\] Control_Unit.C\[19\] Control_Unit.Q\[19\] _0767_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2629_ net5 _1957_ _1896_ net4 _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4315__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4287__I _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4079__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3826__A1 Control_Unit.Q\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4251__A1 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2565__A1 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2868__A2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4490__A1 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2445__I Control_Unit.cont\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2980_ _2304_ _2306_ _2307_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4242__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3596__A3 Control_Unit.Q\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ _0341_ _1655_ _1656_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3601_ _0683_ _0686_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput10 n[2] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4581_ _1985_ _1436_ _1598_ _1602_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3532_ Control_Unit.T\[8\] _2001_ Control_Unit.Q\[8\] _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3463_ _0543_ _0547_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2414_ Control_Unit.cont\[12\] _1724_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3394_ Control_Unit.Rcont _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2345_ Control_Unit.presente\[0\] _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4015_ _1776_ Control_Unit.Q\[9\] _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4481__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4233__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3587__A3 Control_Unit.Q\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4779_ _0103_ net106 Control_Unit.Q\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3511__A3 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2786__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2786__B2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3096__I Control_Unit.T\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2561__I1 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4685__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3018__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2963_ _2280_ _2281_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4702_ _0037_ net57 Control_Unit.cont\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2894_ _1853_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4518__A2 Control_Unit.C\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2529__A1 Control_Unit.cont\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ _1639_ _1641_ _1643_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4564_ _1575_ _1578_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3515_ _0599_ _0614_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout92_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4495_ _1524_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3446_ _0535_ _0550_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3377_ _0497_ _0499_ _0501_ _0502_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4206__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3009__A2 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3248__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__A2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3300_ _0436_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2931__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4280_ _1111_ _1326_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3231_ _0364_ _0365_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3162_ _0237_ _0243_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3093_ _1767_ Control_Unit.T\[8\] _2111_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_35_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3995_ _1776_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _1822_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2877_ _2040_ _2203_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4616_ _1997_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4700__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4547_ _1569_ _1572_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4478_ _0319_ _1491_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3429_ Control_Unit.T\[1\] _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4427__A1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2718__I _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4723__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2800_ _2127_ _2128_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3780_ _0474_ _1976_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2731_ _2059_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ _1990_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4401_ _1418_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3284__I _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2593_ _1809_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4332_ _1915_ Control_Unit.C\[3\] _1802_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4263_ _1286_ _1279_ _1312_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3214_ _0321_ _0325_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4657__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4194_ _1237_ _1235_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3145_ _1821_ _0272_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4409__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3076_ _0214_ _0219_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout55_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3978_ _0238_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2363__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2929_ _1834_ _1944_ _2256_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3148__A1 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3699__A2 Control_Unit.C\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3194__I Control_Unit.Rc vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3320__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2434__I0 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3139__A1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A1 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 n[15] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3862__A2 Control_Unit.Mq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3901_ _0970_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3832_ _0529_ _0901_ _0910_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3763_ _0839_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2714_ _1875_ _2040_ _2042_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3694_ _0767_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2645_ _1705_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2576_ _1903_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3550__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4315_ Control_Unit.C\[1\] _0282_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4246_ _1287_ _1294_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4177_ _1235_ _1233_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2358__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4769__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3128_ _1798_ _0270_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3059_ _1703_ _1687_ _1702_ _0152_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3541__A1 Control_Unit.T\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2731__I _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2430_ _1714_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout105_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2361_ _1689_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4100_ _2037_ _1161_ _1162_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ _1081_ _1083_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3835__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3599__A1 Control_Unit.Q\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4260__A2 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4795_ _0119_ net72 Control_Unit.C\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3815_ Control_Unit.Q\[27\] _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2641__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3746_ _0826_ _0829_ _0830_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3677_ net29 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2628_ _1872_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2559_ net6 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4229_ _0797_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2816__I _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2551__I _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3382__I _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3514__A1 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3817__A2 Control_Unit.C\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2726__I _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3202__B1 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3600_ _0691_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4580_ _1985_ _1601_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput11 n[3] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2556__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3753__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3531_ _0627_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3462_ _0543_ _0547_ _0561_ _0566_ _0553_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_6_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2413_ _1713_ _1723_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3393_ _0510_ _2061_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3505__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2344_ Control_Unit.presente\[2\] _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4014_ _1784_ _1055_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4072__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3992__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2371__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _0102_ net107 Control_Unit.Q\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3729_ Control_Unit.T\[21\] _1981_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2546__I _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4224__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3432__B1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2786__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4160__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2456__I _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4671__I _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2962_ _2280_ _2281_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _0036_ net57 Control_Unit.cont\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3974__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2893_ _1749_ _1754_ _1853_ _2051_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4632_ _0536_ _1642_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3726__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4563_ _1585_ _1586_ _1579_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4494_ _1518_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3514_ _0246_ _2011_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3445_ _0549_ _0278_ _0537_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout85_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3376_ _0497_ _0499_ _0442_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3750__I _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2366__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3197__I _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3925__I _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4142__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3230_ _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2695__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3161_ _0261_ _0269_ _0301_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4436__A2 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3092_ _0235_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3994_ Control_Unit.cont\[5\] Control_Unit.Q\[8\] _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2945_ _2247_ _2259_ _2264_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2876_ _2201_ _2202_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_15_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4615_ _1627_ _1357_ _1624_ _1629_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4546_ _1565_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4477_ _1879_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2922__A2 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__A1 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3428_ _2014_ _0526_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3480__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3359_ _0477_ _0484_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4427__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2824__I _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3938__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2610__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4675__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2913__A2 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A2 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2730_ _1757_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2601__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2661_ Control_Unit.C\[19\] _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4400_ _1356_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3565__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3157__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2592_ _1814_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4331_ _2015_ _1354_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4106__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4262_ _0822_ _0841_ _1299_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3213_ _0348_ _0337_ _0355_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4193_ Control_Unit.Q\[18\] _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3144_ _0281_ _0286_ _0287_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4409__A2 Control_Unit.C\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3075_ _0215_ _0217_ _0218_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2683__A4 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3093__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2840__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2840__B2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3977_ _1040_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2928_ _2255_ _1834_ _1917_ _1911_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4698__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2859_ _1974_ _1975_ _2025_ _2187_ Control_Unit.futuro\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4345__A1 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4529_ _1542_ _1462_ _1554_ _1556_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_2_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3084__A1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2831__A1 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2434__I1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3139__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2898__A1 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4639__A2 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3334__B _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3847__B1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 n[1] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_18_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3075__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2464__I _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3900_ _0971_ _0955_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3831_ _0906_ _0908_ _0909_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3762_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2713_ _2041_ _2040_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3693_ _0771_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2644_ _1676_ _1678_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2889__A1 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2575_ _1762_ _1718_ _1778_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4245_ _0814_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4176_ _1225_ _1227_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3127_ _1799_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3058_ _0197_ _0198_ _0202_ _0203_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2374__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2813__A1 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3541__A2 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__B1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3780__A2 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ net15 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3532__A2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4030_ _1049_ _1070_ _1071_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_38_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4548__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4623__B Control_Unit.C\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4794_ _0118_ net72 Control_Unit.C\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3814_ _0486_ Control_Unit.C\[28\] Control_Unit.Q\[28\] _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3745_ _0826_ _0829_ _0776_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3771__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3676_ _0518_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2627_ _1745_ _1871_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2558_ _1733_ _1886_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4736__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2369__I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2489_ _1809_ _1814_ _1816_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2582__I0 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4228_ _0383_ _0768_ Control_Unit.Q\[19\] _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4159_ Control_Unit.cont\[13\] Control_Unit.Q\[16\] _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3054__A4 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3211__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3514__A2 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3278__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3450__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3450__B2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 n[4] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3059__B _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3530_ _0618_ _0628_ _0626_ _0607_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__4759__CLK net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3461_ _0562_ _0564_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2412_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3392_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2343_ _1676_ _1679_ _1675_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _1838_ _1062_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3748__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3441__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3992__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4777_ _0101_ net107 Control_Unit.Q\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3728_ Control_Unit.Q\[21\] _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3659_ _0734_ _0739_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3483__I Control_Unit.Q\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3432__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3499__A1 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2961_ _1780_ _2231_ _2233_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4700_ _0035_ net59 Control_Unit.cont\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2472__I _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2892_ _2218_ _2219_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _0375_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4562_ _1550_ _1567_ _1568_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2529__A3 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4493_ _1520_ _1522_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3513_ _0246_ _2011_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3444_ _0549_ _0278_ _0537_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3375_ _0500_ _0459_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout78_I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3662__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2382__I Control_Unit.cont\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2940__A3 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3405__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3160_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3091_ _0230_ _0234_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2695__A2 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2416__B _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3993_ _1831_ _1043_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2944_ _2267_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2875_ _2201_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _1353_ _1628_ _1627_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4545_ _1708_ _1988_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4476_ _2036_ Control_Unit.C\[13\] _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3427_ _0531_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3358_ Control_Unit.T\[28\] _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2377__I Control_Unit.cont\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3289_ Control_Unit.T\[18\] _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input10_I n[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4060__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2913__A3 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3874__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4007__I Control_Unit.Q\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2601__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ Control_Unit.C\[16\] _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2591_ _1799_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4330_ _1357_ _1369_ _1371_ _1365_ _0541_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _1286_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3212_ _0350_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4192_ _0996_ _1249_ _1250_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input2_I n[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3143_ _0283_ _0285_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3074_ _2055_ _0216_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4290__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ _1848_ _1042_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2927_ _1825_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2660__I Control_Unit.C\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2858_ _1702_ _2185_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2789_ _2051_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4528_ _1514_ _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4459_ _2046_ Control_Unit.C\[12\] _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4536__B _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2831__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3139__A3 Control_Unit.T\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4336__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3847__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3847__B2 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3350__B _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3830_ _0906_ _0908_ _0522_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3761_ _0840_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2712_ _1711_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3692_ _0754_ _0757_ _0763_ _0772_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_9_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2643_ _1965_ _1969_ _1971_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2574_ _1849_ _1847_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _1348_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4244_ _1283_ _1285_ _1293_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4175_ _0939_ _1232_ _1233_ _0936_ _1234_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout60_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3126_ Control_Unit.T\[3\] _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3057_ _1682_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3066__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2813__A2 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A1 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2577__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3959_ _1025_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4318__A2 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3541__A3 Control_Unit.Q\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2568__A1 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2740__A1 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3532__A3 Control_Unit.Q\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4688__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3048__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4245__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3813_ _0889_ _0892_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4793_ _0117_ net64 Control_Unit.C\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3744_ _0812_ _0827_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3675_ _0725_ _0753_ _0727_ _0764_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2626_ net4 _1896_ _1897_ _1696_ _1954_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3508__B1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _1739_ _1885_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2488_ _1801_ _1811_ _1796_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2582__I1 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4227_ _0788_ _1267_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4158_ _1712_ _1204_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2385__I Control_Unit.cont\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _1139_ _1134_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_3_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3109_ Control_Unit.T\[5\] _2255_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__A1 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3278__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 n[5] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout110_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2961__A1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3460_ _0563_ _0558_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2411_ _1726_ _1738_ _1739_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3391_ _0509_ _1844_ _1842_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2713__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2342_ _1678_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3269__A2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4012_ _1077_ _1063_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4776_ _0100_ net107 Control_Unit.Q\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3727_ _0447_ Control_Unit.C\[22\] Control_Unit.Q\[22\] _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_14_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2952__A1 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3658_ _0735_ _0738_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2952__B2 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3589_ Control_Unit.T\[11\] _2002_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2609_ _1937_ _1932_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3680__A2 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4710__D _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2943__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4448__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3120__A1 _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3671__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2753__I _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2960_ _2283_ _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__B1 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2891_ _2217_ _2211_ _2213_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_30_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4630_ _0281_ _1640_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4561_ _1991_ _1572_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2934__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4492_ _0322_ _1503_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3512_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3443_ _0531_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ Control_Unit.T\[30\] _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3111__A1 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4611__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4759_ _0083_ net55 Control_Unit.Q\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2925__A1 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3350__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2392__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3090_ _2060_ _0232_ _0233_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2695__A3 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3644__A2 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2483__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3992_ _1824_ _0611_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2943_ _2133_ _2257_ _2270_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_15_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2874_ _2045_ _1890_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4613_ _1620_ _1623_ _1356_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4544_ _2176_ _1989_ _1559_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _1492_ _1494_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout90_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3426_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3357_ _0485_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3288_ _0416_ _0396_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2393__I _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3399__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3626__A2 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4051__A2 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2590_ _1913_ _1916_ _1918_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ _0822_ _0841_ _1294_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4191_ _0743_ _1014_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3211_ _0351_ _0352_ _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2478__I _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3142_ _0283_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3073_ _2055_ _0216_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3617__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3093__A3 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4042__A2 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3975_ _1783_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2926_ _2251_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2857_ _1680_ _1685_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2788_ _2069_ _2081_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3553__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4527_ _1544_ _1553_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4458_ _1482_ _1484_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3409_ net19 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4389_ _1425_ _1423_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3608__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3544__A1 Control_Unit.Q\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3760_ _0841_ _0842_ _0843_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2711_ _1860_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3691_ net31 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2642_ _1731_ _1885_ _1887_ _1970_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_12_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2573_ _1764_ _1850_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3535__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _1350_ _1351_ _1355_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4243_ _0822_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4174_ Control_Unit.Q\[16\] _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3125_ _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3056_ _0199_ _0200_ _0201_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout53_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4263__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4015__A2 Control_Unit.Q\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2671__I Control_Unit.C\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2577__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3958_ _0245_ _1026_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2909_ _2227_ _2230_ _2236_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3889_ _0542_ _0951_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3462__B1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3677__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4713__D _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3517__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2740__A2 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3812_ _0876_ _0879_ _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2491__I _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4792_ _0116_ net63 Control_Unit.C\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3756__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3743_ _0813_ _0817_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3674_ _0758_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _1901_ _1952_ _1953_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3508__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4181__A1 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2556_ _1741_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2487_ _1815_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _1194_ _1229_ _1281_ _1230_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4157_ _1736_ _0714_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4484__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3108_ _2067_ _0248_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _1149_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3039_ _1690_ _0160_ _0162_ _0184_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3995__A1 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4782__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2798__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3747__A1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4708__D _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4227__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3986__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3200__I _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3738__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2410__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3202__A3 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 n[6] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4163__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2410_ _1734_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3390_ _0508_ _2068_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2713__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2341_ _1673_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3870__I Control_Unit.Mq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3910__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ _1766_ _1064_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4218__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3311__S _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3110__I Control_Unit.T\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4775_ _0099_ net106 Control_Unit.Q\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2401__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3726_ _0807_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3657_ _0744_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3588_ Control_Unit.T\[11\] _2002_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2608_ net10 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2539_ Control_Unit.cont\[11\] _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4209_ _1261_ _1259_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3968__A1 _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4393__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4678__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2943__A2 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4145__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3904__B _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2459__A1 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3120__A2 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2890_ _2211_ _2213_ _2217_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4560_ _1983_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3865__I _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4491_ _1880_ _1507_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3511_ Control_Unit.T\[7\] Control_Unit.C\[7\] _0611_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3442_ _0543_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_13_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3373_ _0468_ _0469_ _0491_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3111__A2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4827_ _0151_ net89 Control_Unit.T\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4375__A1 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4758_ _0082_ net55 Control_Unit.Q\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3709_ Control_Unit.T\[21\] Control_Unit.C\[21\] Control_Unit.Q\[21\] _0796_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4689_ _0024_ net96 Control_Unit.T\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4127__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3653__A3 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2861__A1 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4602__A2 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4366__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4118__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2392__A3 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3991_ _1839_ _1057_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2942_ _2268_ _2256_ _2269_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2873_ _1745_ _1863_ _1744_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4612_ _1995_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4543_ _1566_ _1567_ _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2907__A2 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4474_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3425_ _0278_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3356_ _0483_ _0480_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3287_ _0409_ _0419_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2674__I _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3399__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3719__B _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2834__A1 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3011__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3562__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4190_ _1236_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3210_ _0317_ _0318_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4511__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3141_ _1925_ _0279_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3072_ Control_Unit.T\[10\] _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2825__A1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ _1773_ Control_Unit.Q\[7\] _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3250__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2925_ _2145_ _2252_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2856_ _2169_ _2181_ _2182_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2787_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4526_ _1544_ _1553_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3553__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4457_ _1480_ _1485_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3408_ _0516_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4388_ _1411_ _1417_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3339_ _0380_ _0470_ _0464_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3963__I _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2710_ _2038_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3690_ _0765_ _0766_ _0778_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2641_ net8 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2572_ _1697_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4311_ _0525_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4242_ _0940_ _1295_ _1296_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _1228_ _1231_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3124_ _0266_ _0267_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3055_ _2190_ _2193_ _2196_ _2206_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_36_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3957_ _1002_ _1008_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2908_ _2061_ _2234_ _2235_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3888_ _0947_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2839_ _2163_ _2166_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2901__B _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2399__I Control_Unit.cont\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4509_ _1530_ _1527_ _1537_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3462__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3453__A1 Control_Unit.C\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3811_ _0868_ _0887_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _0115_ net63 Control_Unit.C\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3742_ _0818_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3673_ _0759_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2624_ net3 _1897_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2555_ _1872_ _1878_ _1744_ _1883_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2486_ _1795_ _1800_ _1810_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4225_ _1280_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4156_ _0996_ _1215_ _1216_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3692__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3107_ _0247_ _0249_ _0250_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4087_ _0317_ _1127_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3038_ _2123_ _0161_ _0171_ _0183_ _0166_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2682__I Control_Unit.C\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4172__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2486__A2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2592__I _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3738__A2 Control_Unit.C\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput15 n[7] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2961__A3 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2340_ Control_Unit.presente\[1\] _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4010_ _1061_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3729__A2 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _0098_ net114 Control_Unit.Q\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3725_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3656_ Control_Unit.Q\[16\] _0745_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3587_ _0345_ Control_Unit.C\[12\] Control_Unit.Q\[12\] _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2607_ net10 _1932_ _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2538_ _1851_ _1855_ _1861_ _1866_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4809__D _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4208_ _1251_ _1115_ _1264_ _1265_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2469_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4139_ _1184_ _1186_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4393__A2 Control_Unit.C\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2587__I _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3656__A1 Control_Unit.Q\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4081__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__A2 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2395__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3510_ Control_Unit.Q\[7\] _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ _2026_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3441_ _0544_ _0545_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4772__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3372_ _0486_ _0495_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__I _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3830__B _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4217__I _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4826_ _0150_ net81 Control_Unit.T\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4757_ _0081_ net53 Control_Unit.Q\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3708_ net32 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4688_ _0023_ net97 Control_Unit.T\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3639_ _0715_ _0729_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2861__A2 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2356__B _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4063__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2613__A2 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4795__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3877__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4054__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3990_ _1042_ _1044_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3876__I _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2941_ _1833_ _1943_ _1835_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2872_ _2045_ _2192_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _1407_ _1625_ _1626_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4542_ _1546_ _1547_ _1545_ _1559_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4473_ _1490_ _1495_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3424_ Control_Unit.Q\[0\] _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3868__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3355_ Control_Unit.T\[27\] _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout76_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2540__A1 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3286_ Control_Unit.T\[17\] _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4809_ _0133_ net106 Control_Unit.C\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3859__B2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3859__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4036__A1 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2365__A4 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3140_ _1812_ Control_Unit.T\[1\] _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3071_ _1857_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4275__A1 Control_Unit.Q\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2825__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3973_ _1825_ _1021_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2924_ _1917_ _1911_ _2249_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2855_ _1967_ _2174_ _2183_ _1725_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_31_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4525_ _1551_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2786_ net17 _2110_ _2114_ net16 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_8_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _2003_ _1462_ _1487_ _1488_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3407_ Control_Unit.Rcont _1730_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4387_ _1405_ _1407_ _1419_ _1424_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _0468_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3269_ _0406_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_27_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4018__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2504__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2809__B _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4009__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2640_ _1968_ _1739_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4050__I _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2571_ _1898_ _1899_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2743__A1 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4310_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4241_ _0814_ _1274_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4172_ _1228_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3123_ _0245_ _0253_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3054_ _1889_ _1737_ _2183_ _2197_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3471__A2 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4225__I _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4420__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3956_ _1002_ _1008_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2907_ _2232_ _2233_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_17_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3887_ _0956_ _0959_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2838_ net6 _2102_ _2165_ _1700_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2769_ _2033_ _2092_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4508_ _1531_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4439_ _1472_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4487__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4239__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2501__A4 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3462__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4175__B1 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2725__A1 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2500__I1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__I Control_Unit.Mq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3810_ _0871_ _0863_ _0881_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4790_ _0114_ net63 Control_Unit.C\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3741_ _0821_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2964__A1 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3756__A3 Control_Unit.Q\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3672_ _0743_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2623_ net17 _1900_ _1902_ _1698_ _1951_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2554_ _1882_ _1877_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2485_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ _1253_ _1276_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _0714_ _1014_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3692__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3106_ _1848_ Control_Unit.T\[7\] _1767_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4086_ _1120_ _1126_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3444__A2 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3037_ _0181_ _0182_ _0170_ _1693_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_24_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3939_ _0990_ _0992_ _0989_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3132__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2486__A3 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 n[8] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3123__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2783__I _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4623__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4773_ _0097_ net114 Control_Unit.Q\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3724_ _0802_ _0808_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _0403_ _1989_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2606_ _1934_ _1928_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3119__I _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3586_ _0676_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2537_ _1862_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2468_ _1796_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4207_ _1254_ _1263_ _1136_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2399_ Control_Unit.cont\[15\] _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4138_ _1184_ _1186_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4069_ _1116_ _1117_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_28_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A1 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2928__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3473__B _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3105__A1 _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__A1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4081__A2 Control_Unit.Q\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2919__A1 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2395__A2 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3440_ _2013_ _0536_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3371_ Control_Unit.T\[30\] _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3647__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4825_ _0149_ net69 Control_Unit.T\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ _0080_ net80 Control_Unit.Q\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3707_ _0725_ _0779_ _0727_ _0794_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4687_ _0022_ net105 Control_Unit.T\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3638_ _0715_ _0729_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3293__B _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3569_ Control_Unit.T\[10\] Control_Unit.C\[10\] _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3312__I _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2598__I _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3877__A2 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2940_ _1788_ _1794_ _2265_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2871_ _2197_ _2198_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _1514_ _1623_ _1620_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4541_ _1562_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4472_ _2018_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3317__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3423_ net30 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3868__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3354_ _0377_ _0479_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2540__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3285_ _0414_ _0415_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout69_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4808_ _0132_ net98 Control_Unit.C\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4739_ _0063_ net101 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3308__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4762__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3070_ _2208_ _0213_ _2037_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3972_ _1819_ _0599_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2923_ _2249_ _2250_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2854_ _2177_ _1967_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2785_ _2113_ _2083_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4524_ _1533_ _1535_ _1549_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4455_ _1479_ _1486_ _1421_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3406_ _0515_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4386_ _1422_ _1423_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3337_ _0463_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3268_ _0388_ _0398_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3199_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4785__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4018__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout119_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2570_ _1748_ _1753_ _1853_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _1292_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4171_ _1194_ _1229_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3122_ _0263_ _1916_ _0265_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4248__A2 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3053_ _2199_ _2311_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3471__A3 Control_Unit.Q\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3410__I Control_Unit.Mx vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3955_ _2067_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2906_ _2232_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4420__A2 Control_Unit.C\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3886_ _0956_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4184__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2837_ _1700_ _2165_ _2107_ _1695_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2768_ _2029_ _2094_ _2096_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2699_ _2027_ _1876_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4507_ _1533_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3931__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _1466_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2498__A1 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4369_ _1406_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4175__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2725__A2 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2489__B2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2489__A1 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2555__B _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2413__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3740_ _0822_ _0823_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ Control_Unit.T\[17\] _1987_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2622_ _1906_ _1949_ _1950_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2553_ _1881_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3913__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2484_ _1812_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4223_ _1266_ _1270_ _1277_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4154_ _1212_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4085_ _0351_ _1148_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3105_ _0239_ _0248_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3036_ _1929_ _1931_ _0173_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3444__A3 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2465__B _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4823__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3938_ _2070_ _1002_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3869_ _0506_ _0531_ _0943_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4157__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3380__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4632__A2 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2375__B _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2643__A1 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput17 n[9] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4148__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4320__A1 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4387__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4772_ _0096_ net114 Control_Unit.Q\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3723_ _0796_ _0800_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3654_ _0403_ Control_Unit.C\[16\] _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2605_ _1933_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3585_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2536_ _1863_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout99_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2467_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4206_ _1254_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4311__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2398_ _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4137_ _2177_ _1188_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2873__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3019_ _2254_ _2258_ _0164_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_36_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4378__A1 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4719__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4302__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2616__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4604__I _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2919__A2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3370_ _0495_ _0494_ _0489_ _0496_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_fanout101_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2794__I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2607__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4824_ _0148_ net64 Control_Unit.T\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4755_ _0079_ net53 Control_Unit.Q\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3706_ _0786_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4686_ _0021_ net106 Control_Unit.T\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3637_ _0718_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4532__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3568_ Control_Unit.T\[10\] Control_Unit.C\[10\] _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2519_ _1717_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3499_ _0254_ _2007_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3099__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4048__B1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3023__A1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4691__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2837__B2 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2837__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3262__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2870_ _2190_ _2193_ _2196_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_43_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _1544_ _1553_ _1551_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4471_ _1349_ _1497_ _1501_ _1365_ _1502_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2789__I _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3422_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3868__A3 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3353_ _0482_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3284_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4293__A3 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _0131_ net100 Control_Unit.C\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2999_ _2277_ _2278_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4738_ _0062_ net97 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4669_ _1668_ _1670_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4505__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4275__A3 Control_Unit.Q\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ _2070_ _1038_ _1039_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2922_ _1918_ _1829_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3786__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2853_ _1970_ _2097_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2784_ _2112_ _1780_ _2062_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4499__B1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4454_ _1479_ _1486_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3405_ _0511_ _2174_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4385_ _1410_ _1418_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3344__S _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3336_ _0400_ _0401_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout81_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3267_ _1966_ _0386_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3198_ Control_Unit.Mt _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3226__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3529__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3701__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3988__I _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3768__A2 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2991__A3 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4612__I _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2743__A3 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4170_ _1211_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3121_ _1826_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3052_ _1970_ _2313_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3456__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4653__B1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3759__A2 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ _1018_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2905_ _1781_ _1899_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3885_ _0958_ _0948_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2836_ _2164_ _2089_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2767_ _1730_ _1874_ _2095_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2698_ _2026_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4506_ _1707_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _1468_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4368_ Control_Unit.Mc _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3319_ _0448_ _0450_ _0451_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _0927_ _1274_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2670__A2 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2973__A3 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3492__B _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2489__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4754__D _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__I _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2413__A2 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3670_ Control_Unit.T\[17\] _1987_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2621_ net16 _1902_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2552_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4775__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4222_ _1261_ _1269_ _1259_ _1245_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2483_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4153_ _1213_ _1194_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4084_ _1142_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3104_ _2070_ _0246_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3035_ _0180_ _0174_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3421__I Control_Unit.Mx vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3937_ _0979_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3601__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3868_ _0282_ _1804_ _0544_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4157__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2819_ _2147_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3799_ _0876_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3668__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2375__C _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 start net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4798__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4320__A2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3241__I _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2634__A2 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _0095_ net112 Control_Unit.Q\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4387__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3722_ _0796_ _0800_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3653_ _0413_ Control_Unit.C\[17\] _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2604_ _1797_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3584_ _0670_ _0678_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2535_ Control_Unit.cont\[9\] _1747_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2570__A1 _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3416__I _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2466_ Control_Unit.cont\[2\] _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4205_ _1259_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4311__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ _1182_ _1187_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2397_ _1710_ _1725_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2873__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ _1128_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3018_ _2263_ _2275_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4378__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3050__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3889__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3326__I _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4066__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3813__A1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2616__A2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3236__I _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4813__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4057__A1 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4823_ _0147_ net81 Control_Unit.T\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4754_ _0078_ net53 Control_Unit.Q\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3705_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4685_ _0020_ net98 Control_Unit.T\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3636_ _0701_ _0705_ _0711_ _0719_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4532__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3567_ Control_Unit.T\[11\] _2002_ Control_Unit.Q\[11\] _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3146__I Control_Unit.T\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2543__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ _1830_ _1837_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3498_ _0598_ Control_Unit.C\[6\] _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2449_ _1761_ _1777_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_5_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4119_ _1165_ _1167_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4048__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3271__A2 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3023__A2 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3262__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4211__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _2019_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3421_ Control_Unit.Mx _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2525__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3352_ _0480_ _0481_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3283_ Control_Unit.Rc _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4450__A1 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3253__A2 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3789__B1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _0130_ net99 Control_Unit.C\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2998_ _2247_ _2259_ _2264_ _2272_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4737_ _0061_ net85 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4668_ _0313_ _1640_ _1669_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4505__A2 Control_Unit.C\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3619_ _0623_ _0700_ _0625_ _0712_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4599_ _1612_ _1613_ _1979_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4441__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2755__A1 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2755__B2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2507__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3180__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4757__D _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3970_ _1020_ _1022_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2921_ _1821_ _1917_ _1805_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2852_ _2172_ _2175_ _2180_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_31_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2783_ _2111_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _1533_ _1535_ _1549_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2746__A1 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4453_ _1480_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3404_ _0514_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4499__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4384_ _1421_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2749__B _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3335_ _0425_ _0461_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout74_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3266_ _0404_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3197_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3226__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4423__A1 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2503__I _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2976__A1 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3509__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2900__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ _0262_ _2073_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3051_ _1970_ _2313_ _2314_ _1964_ _0196_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3953_ _1783_ _1020_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2904_ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3884_ _1926_ _0953_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2835_ _2054_ _2088_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2719__A1 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2766_ _1966_ _1874_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2697_ _1734_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4505_ _1879_ Control_Unit.C\[15\] _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ _0238_ _2000_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3144__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4367_ _2011_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3318_ Control_Unit.T\[20\] _0445_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_24_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _1033_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3249_ _1882_ _0366_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2670__A3 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2958__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3135__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2949__B2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2949__A1 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3239__I _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2620_ _1689_ _1905_ _1908_ _1691_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2551_ _1879_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2482_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4221_ _1247_ _1252_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4323__B1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4152_ _1189_ _1191_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4083_ _0322_ _1144_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_37_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3103_ _0245_ _0246_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4626__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3034_ _2274_ _2141_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3936_ _1004_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3867_ _0549_ _0937_ _0940_ _0942_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2818_ _1688_ _2145_ _2142_ _1937_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3798_ Control_Unit.Q\[26\] _0877_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3365__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2749_ _2074_ _2076_ _2072_ _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3668__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4419_ _1441_ _1450_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__A2 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3108__A1 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _0094_ net112 Control_Unit.Q\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ _0780_ _0785_ _0793_ _0801_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_14_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3652_ Control_Unit.Q\[17\] _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3583_ _0664_ _0677_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2603_ _1929_ _1930_ _1931_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2534_ Control_Unit.cont\[10\] _1858_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2570__A2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2465_ _1789_ _1790_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4204_ _1261_ _1245_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2396_ _1711_ _1712_ _1724_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_25_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ _1177_ _1115_ _1194_ _1196_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4066_ _0222_ _1129_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3017_ _1690_ _0160_ _0162_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3919_ _0967_ _0969_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3338__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3889__A2 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4765__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3813__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3329__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3501__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _0146_ net69 Control_Unit.T\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4753_ _0077_ net55 Control_Unit.Q\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3704_ _0787_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4684_ _0019_ net98 Control_Unit.T\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ _0523_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ net21 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3740__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2517_ _1840_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3497_ Control_Unit.Q\[6\] _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2448_ _1772_ _1775_ _1776_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2379_ _1707_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4118_ _1165_ _1167_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4049_ Control_Unit.Q\[11\] _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input17_I n[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4207__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3559__A1 Control_Unit.T\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2950__B _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3337__I _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3731__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3798__A1 Control_Unit.Q\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4631__I _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3247__I _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3420_ _0517_ _0519_ _0524_ _0527_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3351_ _0380_ _0470_ _0476_ _0478_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3282_ _0413_ _0363_ _0341_ _0420_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I n[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3238__B1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3789__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4805_ _0129_ net114 Control_Unit.C\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2997_ _1697_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4736_ _0060_ net96 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2764__A2 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4667_ _0235_ _0332_ _0333_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3618_ _0706_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3713__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _0490_ _1615_ _1353_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3549_ _0644_ _0646_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2755__A2 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3180__A2 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2920_ _1916_ _1933_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4196__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2851_ _2172_ _2179_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4196__B2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2782_ _1759_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4521_ _1545_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2746__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4452_ _1482_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3403_ _0511_ _2173_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4383_ _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3334_ _0422_ _0465_ _0342_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3265_ _0384_ _0403_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_6_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout67_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3196_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4423__A2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ Control_Unit.futuro\[2\] net71 Control_Unit.presente\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A2 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output48_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2728__A2 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3525__I _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3050_ _1888_ _2317_ _0195_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4102__A1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4653__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2416__A1 _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ _1785_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2903_ _1764_ _2061_ _1854_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3883_ _1813_ _0544_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2834_ _1695_ _2107_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2604__I _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3916__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _0351_ _1528_ _1532_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2765_ _2031_ _2032_ _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2696_ _1680_ _1674_ _1683_ _2024_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4435_ _1852_ _1455_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3435__I Control_Unit.C\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4366_ _1350_ _1402_ _1404_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3317_ _0430_ _0435_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ _0927_ _1334_ _1341_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3248_ _1882_ _0366_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3179_ _0222_ _0213_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4644__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4580__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3135__A2 Control_Unit.T\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4332__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4635__A2 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4399__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2949__A2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__B _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2550_ _1712_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout117_I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2481_ _1770_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4220_ _1263_ _1270_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4323__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4151_ _1210_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2885__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _2046_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3102_ Control_Unit.T\[6\] _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3033_ _1698_ _2333_ _0160_ _1690_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_37_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3935_ _1914_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3866_ _0941_ _0549_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2817_ _1688_ _2145_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3797_ _0477_ Control_Unit.C\[26\] _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2748_ _1793_ _1918_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4418_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2679_ Control_Unit.C\[4\] _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _1367_ _1373_ _1376_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2628__A1 _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2509__I _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2867__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4634__I _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3044__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3720_ net33 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3651_ net27 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4544__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3582_ _0664_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2602_ _1927_ net9 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2533_ _1716_ _1748_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2464_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4203_ _1239_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2395_ _1713_ _1723_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2858__A1 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4134_ _1192_ _1195_ _0976_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4065_ _1098_ _1103_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3016_ _2123_ _0161_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3918_ _1926_ _0965_ _0966_ _0969_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_20_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3849_ _0925_ _0923_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2849__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4471__B1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__I _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3265__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _0145_ net68 Control_Unit.T\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3568__A2 Control_Unit.C\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4752_ _0076_ net77 Control_Unit.Q\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3703_ _0788_ _0789_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4683_ _0018_ net111 Control_Unit.T\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4517__A1 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3634_ net26 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3565_ _0518_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2516_ _1761_ _1777_ _1842_ _1844_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout97_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3496_ Control_Unit.T\[6\] _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4539__I _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2447_ Control_Unit.cont\[6\] _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3443__I _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2378_ _1706_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4117_ _1174_ _1171_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4048_ _1056_ _1109_ _1110_ _1112_ _1113_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3008__A1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3559__A2 Control_Unit.C\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2950__C _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4223__B _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3722__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3350_ _0422_ _0479_ _0342_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3281_ _0418_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2461__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4804_ _0128_ net110 Control_Unit.C\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2996_ net4 _2321_ _2323_ _1696_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4735_ _0059_ net85 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3438__I Control_Unit.Q\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4666_ _0216_ _1642_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3617_ _0707_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4597_ _1612_ _1979_ _1608_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4755__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3548_ _0644_ _0646_ _0539_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2921__B1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3173__I _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3479_ _0518_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3477__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3229__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3401__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3348__I _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3704__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2850_ _2174_ _2173_ _2178_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2781_ _2058_ _2084_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_15_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4520_ _1546_ _1547_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4778__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4451_ _2060_ _2004_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3402_ _0513_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4382_ _0421_ _1352_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3333_ _0462_ _0463_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3264_ _0384_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3459__A1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3195_ _0338_ Control_Unit.Mt _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4187__A2 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2979_ _1751_ _2216_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4718_ Control_Unit.futuro\[1\] net57 Control_Unit.presente\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4649_ _0254_ _1642_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2370__A1 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3078__I _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3806__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4350__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ _1769_ Control_Unit.Q\[6\] _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2416__A2 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2902_ _2118_ _2226_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3882_ _1799_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2833_ _2109_ _2160_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2764_ _2033_ _2092_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4503_ _2027_ _1519_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2695_ _1980_ _1999_ _2005_ _2023_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4434_ _2046_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4365_ _2007_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3316_ _0400_ _0401_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _1335_ _1341_ _0927_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3247_ _1710_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3178_ _1713_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4332__A2 Control_Unit.C\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2646__A2 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2480_ _1808_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4150_ _1197_ _1198_ _1209_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3101_ _1832_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4087__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4081_ _1715_ Control_Unit.Q\[12\] _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4367__I _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3032_ _2123_ _0161_ _0166_ _0177_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3934_ _1795_ Control_Unit.Q\[5\] _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3865_ _2153_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2816_ _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4011__A1 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3796_ _0477_ Control_Unit.C\[26\] _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2747_ _1828_ _1806_ _2075_ _2074_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2678_ _2006_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4417_ _1442_ _1449_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_8_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4348_ _1382_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4078__A1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4279_ _1112_ _1326_ _1327_ _1328_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3044__A2 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3650_ _0725_ _0726_ _0727_ _0741_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3581_ _0667_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2601_ _1921_ net2 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2555__A1 _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2532_ _1856_ _1860_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4202_ _1241_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2463_ _1791_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2394_ _1714_ _1715_ _1716_ _1722_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__2858__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4133_ _1178_ _1179_ _1172_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ _1098_ _1103_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3015_ _0156_ _0158_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4560__I _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3917_ _0979_ _0982_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3848_ _0917_ _0920_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3779_ _0474_ Control_Unit.C\[25\] _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2849__A2 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout110 net112 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4470__I _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2785__A1 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2537__A1 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3734__B1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4462__A1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4820_ _0144_ net68 Control_Unit.T\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _0075_ net96 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3702_ Control_Unit.T\[19\] _1990_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4682_ _0017_ net115 Control_Unit.T\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4517__A2 Control_Unit.C\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3633_ _0528_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3564_ _0623_ _0649_ _0625_ _0661_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2515_ _1843_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3495_ net47 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2446_ _1773_ _1774_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2377_ Control_Unit.cont\[15\] _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4116_ _1139_ _1134_ _1152_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_25_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4047_ Control_Unit.Q\[10\] _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4684__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3008__A2 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3707__B1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3280_ _0413_ _0414_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2930__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3238__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4435__A1 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _0127_ net113 Control_Unit.C\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2995_ _2299_ _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4734_ _0058_ net82 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2749__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4665_ _1665_ _1667_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3616_ Control_Unit.Q\[13\] _0708_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4596_ _1612_ _1610_ _1614_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3547_ _0631_ _0636_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2921__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3478_ _0529_ _0574_ _0524_ _0581_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2429_ _1757_ _1722_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3229__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2912__A1 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4114__B1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2708__I _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2979__A1 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2780_ net3 _2108_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2600__B1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4450_ _2047_ _1467_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3401_ _0511_ _1877_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4381_ _1410_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3332_ Control_Unit.T\[24\] _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3263_ Control_Unit.T\[16\] _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3459__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3194_ Control_Unit.Rc _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3449__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2978_ _2214_ _2305_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4722__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3395__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ Control_Unit.futuro\[0\] net58 Control_Unit.presente\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4648_ _1653_ _1654_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4579_ _0421_ _1600_ _1364_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2370__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2528__I _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3622__A2 Control_Unit.C\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3386__A1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3094__I _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2438__I _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ _1819_ _1005_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2901_ _2225_ _2227_ _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3613__A2 Control_Unit.C\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _0953_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ net3 _2108_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2763_ _2035_ _2044_ _2090_ _2091_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _1520_ _1522_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3129__A1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2694_ _2012_ _2017_ _2022_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4433_ _1752_ Control_Unit.C\[10\] _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4364_ _1352_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3315_ _0410_ _0419_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4295_ _1332_ Control_Unit.Q\[29\] _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout72_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3246_ _0384_ _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3301__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3177_ _0317_ _0318_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_27_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__A2 Control_Unit.C\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3907__I _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4332__A3 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4768__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3359__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2721__I _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3100_ _0237_ _0243_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ _2059_ _1114_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3031_ _1693_ _0170_ _0171_ _0176_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3933_ _1797_ _0986_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3864_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2815_ _1808_ _1813_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3795_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2746_ _1934_ _1812_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2677_ Control_Unit.C\[5\] _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3770__A1 Control_Unit.Q\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4416_ _2001_ _1407_ _1436_ _1451_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3522__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4347_ _1383_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4278_ Control_Unit.Q\[26\] _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3229_ _0367_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3825__A2 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4250__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3637__I _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3761__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3513__A1 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3816__A2 Control_Unit.C\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3321__B _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4241__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2600_ _1927_ net9 net2 _1928_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3580_ _0650_ _0654_ _0660_ _0668_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2531_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3752__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _1255_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2462_ _1773_ _1771_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2393_ _1721_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4132_ _1178_ _1179_ _1193_ _1172_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4063_ _0322_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3014_ _2247_ _0159_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_3_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4480__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4232__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3916_ _1915_ _0985_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2361__I _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3847_ _0832_ _0911_ _0834_ _0924_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3991__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3778_ Control_Unit.T\[26\] Control_Unit.C\[26\] Control_Unit.Q\[26\] _0860_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2729_ _2055_ _2056_ _2057_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4299__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout111 net112 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout100 net109 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4806__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2785__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3734__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3734__B2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4462__A2 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4750_ _0074_ net102 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3701_ Control_Unit.T\[19\] _1990_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4681_ _0016_ net111 Control_Unit.T\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3973__A1 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3632_ _0662_ _0713_ _0724_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3563_ _0655_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2514_ _1719_ _1720_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3494_ _0582_ _0583_ _0596_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2445_ Control_Unit.cont\[5\] _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ Control_Unit.Q\[14\] _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2376_ _1704_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4141__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3955__A1 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3707__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3707__B2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3046__B _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2930__A2 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2446__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4199__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4802_ _0126_ net113 Control_Unit.C\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2994_ _2294_ _2298_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4733_ _0057_ net82 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3946__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4664_ _0332_ _1640_ _1666_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3615_ _0349_ _2018_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4595_ _1612_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3546_ _0632_ _0635_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3477_ _0578_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2428_ Control_Unit.cont\[8\] _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3470__I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2359_ net9 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4029_ _1092_ _1087_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input15_I n[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2676__A1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3928__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2600__A1 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2600__B2 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3400_ _0509_ _2191_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4353__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4380_ _1411_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2903__A2 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4674__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3331_ _0448_ _0461_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4105__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3262_ _0400_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3193_ _0220_ _0335_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input7_I n[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A2 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2977_ _2215_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3395__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4716_ _0000_ _4716_/E _4716_/RN Control_Unit.Rcont vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__3465__I _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _0297_ _0268_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4344__A1 Control_Unit.C\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4578_ _1584_ _1592_ _1599_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3529_ _0613_ _0616_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2370__A3 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3083__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3622__A3 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4583__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3386__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2897__A1 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3074__A1 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2900_ _1755_ _2212_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3613__A3 Control_Unit.Q\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _1800_ _1810_ Control_Unit.Q\[2\] _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_16_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2831_ _1697_ _2110_ _2116_ _2152_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2762_ _2034_ _2042_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4501_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2693_ _2018_ _2019_ _2020_ _2021_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4432_ _1456_ _1458_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4363_ _1394_ _1396_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3314_ _0414_ _0415_ _0413_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _1339_ _1337_ _1340_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3245_ _2176_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3176_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout65_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2364__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output46_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3833__I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2590__I0 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3030_ _0172_ _0173_ _0175_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3047__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3598__A2 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3932_ _1801_ Control_Unit.Q\[4\] _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3863_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4613__B _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4547__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2814_ _2141_ _2139_ _2142_ _1937_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3794_ Control_Unit.T\[27\] Control_Unit.C\[27\] Control_Unit.Q\[27\] _0875_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2745_ _2073_ _1805_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2676_ _2000_ _2001_ _2003_ _2004_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4415_ _1441_ _1450_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4346_ _1915_ _1384_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2359__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4277_ _1306_ _1322_ _1317_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3228_ _1889_ _0368_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3159_ _0302_ _0258_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3589__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4250__A3 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3210__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3761__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4735__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3513__A2 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3029__A1 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2530_ _1857_ _1858_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout115_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2461_ _1785_ _1719_ _1784_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4200_ _1256_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2392_ _1717_ _1718_ _1719_ _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4131_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4062_ _1120_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3268__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3013_ _0156_ _0158_ _0154_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4232__A3 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _1933_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3846_ _0922_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3777_ net37 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2728_ _1750_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4758__CLK net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2659_ _1987_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout112 net116 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout101 net105 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4329_ _1370_ _1366_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4471__A3 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2552__I _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3383__I Control_Unit.Rcont vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2727__I _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ Control_Unit.Q\[19\] _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4680_ _0015_ net110 Control_Unit.T\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3631_ _0719_ _0722_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3562_ _0656_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2513_ _1841_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3493_ _0592_ _0594_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2444_ Control_Unit.cont\[4\] _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2375_ _1687_ _1688_ _1702_ _1703_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4114_ _1158_ _1115_ _1056_ _1176_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_29_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2637__I _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4045_ Control_Unit.Mq _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3468__I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3829_ _0893_ _0899_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4248__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2547__I _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3891__A1 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2694__A2 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _0125_ net93 Control_Unit.C\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2993_ _2318_ _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4732_ _0056_ net82 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3946__A2 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4663_ _0244_ _0308_ _0310_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3614_ Control_Unit.T\[13\] _2018_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4594_ _1421_ _1608_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3237__B _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3545_ _0640_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout95_I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3476_ _0570_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4123__A2 Control_Unit.Q\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2427_ _1751_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3882__A1 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2358_ net10 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2367__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4028_ _1074_ _0937_ _1056_ _1094_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4582__I _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2373__A1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4114__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2676__A2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3625__A1 Control_Unit.Q\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2600__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4819__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3330_ _0416_ _0396_ _0425_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3261_ _0382_ _0373_ _0392_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3192_ _0326_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3616__A1 Control_Unit.Q\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3520__B _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2976_ _1863_ _2201_ _2202_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4041__A1 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4715_ _0004_ _4715_/E _4715_/RN net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__2650__I Control_Unit.C\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4646_ _0299_ _1651_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4577_ _1981_ _1985_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3528_ _0613_ _0616_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2370__A4 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3459_ _0563_ _0558_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4280__A1 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__A1 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2560__I _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2594__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3605__B _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3074__A2 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2735__I _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2830_ _2121_ _2158_ _2115_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2761_ _2054_ _2088_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4500_ _1518_ _1523_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2692_ Control_Unit.C\[14\] _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4431_ _1459_ _1464_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4326__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4362_ _1397_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4791__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3313_ Control_Unit.T\[22\] _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4293_ _1332_ _1339_ _0976_ _1335_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3244_ Control_Unit.T\[15\] _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3837__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3175_ _2041_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout58_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4262__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3065__A2 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4014__A1 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2959_ _2285_ _2286_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4629_ _0377_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3056__A2 _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3764__B1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2590__I1 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4492__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2893__C _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3047__A2 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3931_ _1821_ _1000_ _1001_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _0338_ Control_Unit.Mq _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2813_ _1928_ _2133_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3793_ _0873_ _0869_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _1820_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2675_ Control_Unit.C\[10\] _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4414_ _1442_ _1449_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4345_ _2015_ _1807_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4276_ _1316_ _1325_ _0946_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3227_ _0320_ _0349_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3158_ _0251_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4687__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3089_ _1768_ _0231_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3277__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4226__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3029__A2 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4529__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2460_ _1772_ _1775_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4130_ _1189_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2391_ Control_Unit.cont\[4\] Control_Unit.cont\[5\] _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4061_ _1857_ _1122_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_7_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3012_ _2259_ _2264_ _0157_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3914_ _1800_ Control_Unit.Q\[4\] _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3845_ _0913_ _0916_ _0921_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3776_ _0765_ _0848_ _0858_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2727_ _2051_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2658_ Control_Unit.C\[17\] _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2703__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout113 net116 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout102 net104 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_2589_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4328_ Control_Unit.C\[0\] _1814_ _1359_ _1361_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4259_ _1309_ _1310_ _1280_ _1211_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4456__A1 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4208__A1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3498__A2 Control_Unit.C\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3670__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3630_ _0719_ _0722_ _0672_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3561_ Control_Unit.Q\[9\] _0657_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2933__A1 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2512_ _1824_ _1772_ _1774_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4135__B1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3492_ _0592_ _0594_ _0539_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2443_ _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2374_ net11 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4113_ _1173_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4044_ _1088_ _1108_ _1096_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2653__I _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3413__A2 Control_Unit.Mx vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4610__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3828_ _0894_ _0898_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3177__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3759_ Control_Unit.T\[23\] _1984_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2860__B1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3394__I Control_Unit.Rcont vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2915__A1 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__A2 Control_Unit.cont\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2694__A3 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3643__A2 Control_Unit.C\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4800_ _0124_ net92 Control_Unit.C\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2992_ _2229_ _2319_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _0055_ net82 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4662_ _0225_ _1644_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3613_ _0362_ Control_Unit.C\[14\] Control_Unit.Q\[14\] _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_31_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _1976_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3544_ Control_Unit.Q\[8\] _0641_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3475_ _0543_ _0547_ _0548_ _0552_ _0571_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2426_ _1754_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout88_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2357_ _1679_ _1682_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4027_ _1090_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2383__I Control_Unit.cont\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3479__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3398__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3570__A1 Control_Unit.Q\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4259__B _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3322__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2676__A3 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3873__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3389__A1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3561__A1 Control_Unit.Q\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3260_ _0387_ _0391_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3191_ _0328_ _0334_ _0314_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2975_ _2220_ _2302_ _2218_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4714_ _0001_ _4714_/E _4714_/RN Control_Unit.Mx vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_30_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4645_ _1651_ _0347_ _1652_ _0397_ _0263_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4576_ _1982_ _1593_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3527_ _0570_ _0579_ _0605_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3304__A1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3458_ _0557_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2409_ _1735_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2378__I _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3389_ _0508_ _2265_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4593__I _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2594__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3846__A2 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4559__B1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2760_ _2039_ _2043_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2691_ Control_Unit.C\[15\] _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4430_ _1447_ _1452_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3534__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _0979_ _1398_ _1399_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3312_ _0446_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4292_ Control_Unit.Q\[29\] _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3243_ _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3174_ Control_Unit.T\[12\] _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4262__A2 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4565__A3 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2958_ _2068_ _2239_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2576__A2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2889_ _1751_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4628_ _0506_ _0532_ _0280_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4559_ _1349_ _1580_ _1582_ _1406_ _1583_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3764__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput50 net50 X[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3930_ _0985_ _0987_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3861_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3792_ _0864_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2812_ net11 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2743_ _1910_ _1816_ _1817_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3755__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2674_ _2002_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4413_ _1447_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4180__A1 Control_Unit.cont\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4344_ Control_Unit.C\[3\] _1807_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4275_ Control_Unit.Q\[24\] _1322_ Control_Unit.Q\[26\] _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout70_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3226_ _0320_ _0349_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2656__I Control_Unit.C\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2494__B2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2494__A1 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3157_ _0277_ _0296_ _0298_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3088_ _1768_ _0231_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3994__A1 Control_Unit.cont\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4171__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4267__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2788__A2 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3985__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4162__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2390_ Control_Unit.cont\[3\] Control_Unit.cont\[2\] Control_Unit.cont\[1\] Control_Unit.cont\[0\]
+ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3860__I Control_Unit.Mq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4060_ _1123_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2476__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3011_ _1944_ _2276_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3976__A1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3913_ _0282_ _0983_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3844_ _0913_ _0916_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4640__B _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3775_ _0854_ _0856_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2400__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2726_ _2050_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2657_ _1982_ _1983_ _1984_ _1985_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_12_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3900__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout103 net104 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2588_ _1816_ _1817_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout114 net115 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4327_ _1367_ _1368_ _1363_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4258_ _1229_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3209_ _0317_ _0318_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4456__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4189_ _1237_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4208__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3431__A3 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3719__A1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4392__A1 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__A1 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3498__A3 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A1 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2630__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3560_ _0225_ Control_Unit.C\[9\] _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4677__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2511_ _1839_ _1789_ _1790_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3491_ _0578_ _0580_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2442_ _1769_ Control_Unit.cont\[2\] Control_Unit.cont\[1\] _1770_ _1771_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2373_ _1694_ _1699_ _1701_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4112_ _1174_ _1156_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _1088_ _1096_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2621__A1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3827_ _0902_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3758_ Control_Unit.T\[23\] _1984_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4374__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2709_ _2037_ _1749_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3689_ _0772_ _0775_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2860__A1 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2860__B2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2612__B2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4711__D _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4668__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4455__B _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3643__A3 Control_Unit.Q\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2991_ _2225_ _2227_ _2228_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_22_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ _0054_ net79 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4661_ _1662_ _1664_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3612_ _0701_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2906__A2 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4592_ _1606_ _1610_ _1611_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3543_ _0231_ Control_Unit.C\[8\] _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3474_ _0575_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2425_ _1753_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3867__B1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2356_ _1680_ _1676_ _1684_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__B1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4026_ _1091_ _1072_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2664__I _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3398__A2 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3495__I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2373__A3 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3322__A2 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2676__A4 _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3086__A1 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3389__A2 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3190_ _0235_ _0332_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2484__I _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2974_ _2229_ _2237_ _2300_ _2301_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4577__A1 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ _0006_ _4713_/E _4713_/RN Control_Unit.Mt vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _0277_ _0296_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4575_ _1982_ _1596_ _1597_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2355__A3 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3526_ _0604_ _0617_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2659__I _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3457_ _0542_ _0556_ _0560_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2408_ _1736_ _1724_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3388_ _0509_ _1816_ _1817_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2339_ Control_Unit.presente\[0\] _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4009_ _2112_ _1066_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I n[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4568__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3240__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4738__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3543__A2 Control_Unit.C\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3059__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2806__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4559__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3231__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2690_ Control_Unit.C\[12\] _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3863__I _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4360_ _2008_ _0971_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3311_ _0443_ _0444_ _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4291_ _1337_ _1338_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3242_ _1707_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3173_ _2037_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I n[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2957_ _2238_ _2284_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2888_ _2214_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4627_ _0533_ _0363_ _1638_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _1991_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2389__I Control_Unit.cont\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4489_ _2041_ Control_Unit.C\[14\] _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3509_ net48 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3461__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3516__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput51 net51 b vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput40 net40 X[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3632__B _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3858__I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3860_ Control_Unit.Mq _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3791_ _0871_ _0863_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2811_ _1703_ _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2742_ _2070_ _1835_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2673_ Control_Unit.C\[11\] _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4412_ _1444_ _1446_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4343_ _1825_ Control_Unit.C\[4\] _1797_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4274_ _1322_ _1323_ _1324_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3225_ _1881_ _0366_ _2177_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_41_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2494__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3156_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3087_ Control_Unit.T\[8\] _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2672__I Control_Unit.C\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3994__A2 Control_Unit.Q\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3989_ _1042_ _1044_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3717__B _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2847__I _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4548__B _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output44_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4714__D _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3985__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2476__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3010_ _0154_ _0155_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2492__I _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3912_ _1811_ _0557_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3843_ _0917_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3774_ _0854_ _0856_ _0776_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2725_ _2045_ _1751_ _2039_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2656_ Control_Unit.C\[22\] _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4153__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout104 net105 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2587_ _1915_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout115 net116 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3272__B _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4326_ _1359_ _1366_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4257_ _1156_ _1307_ _1192_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2667__I Control_Unit.C\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4188_ _1245_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3208_ _1711_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3664__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3139_ _1933_ _0282_ Control_Unit.T\[2\] _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4392__A2 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4709__D _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3407__A1 Control_Unit.Rcont vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout113_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2394__A1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3490_ _0576_ _0564_ _0575_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2510_ _1838_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4135__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2441_ Control_Unit.cont\[0\] _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2372_ net8 net7 net6 _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_25_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4111_ _1149_ _1151_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4042_ _1104_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3646__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3949__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3826_ Control_Unit.Q\[28\] _0903_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3177__A3 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3757_ Control_Unit.Q\[23\] _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4374__A2 Control_Unit.C\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2708_ _2036_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3688_ _0772_ _0775_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2639_ _1967_ _1729_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4771__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2688__A2 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4309_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2612__A2 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4365__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2990_ _2237_ _2300_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4053__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _0308_ _1640_ _1663_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3611_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4591_ _1603_ _1600_ _1609_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3564__B1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4794__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3542_ Control_Unit.T\[8\] Control_Unit.C\[8\] _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3473_ _0563_ _0558_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2424_ _1752_ _1722_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2355_ _1675_ _1679_ _1682_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3619__B2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4025_ _1067_ _1069_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2680__I _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3809_ _0835_ _0838_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4789_ _0113_ net63 Control_Unit.C\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4400__I _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2530__A1 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3086__A2 Control_Unit.T\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2833__A2 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4035__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4310__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2521__A1 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2973_ _2225_ _2227_ _2228_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4577__A2 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4712_ _0003_ _4712_/E _4712_/RN Control_Unit.Mq vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4329__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _0277_ _0296_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4574_ _1982_ _1594_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3525_ _0523_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout93_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3456_ _0542_ _0556_ _0559_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2407_ Control_Unit.cont\[12\] _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3387_ _0507_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2512__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2338_ _1675_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2675__I Control_Unit.C\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4008_ _1059_ _1065_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4265__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4568__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3240__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3059__A2 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2806__A2 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3310_ Control_Unit.T\[21\] _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2742__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4290_ _0947_ _1335_ _1332_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3241_ _0381_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3172_ _0229_ _0313_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2956_ _2064_ _1904_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2887_ _1745_ _1860_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _0506_ _0532_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4557_ _1993_ _1570_ _1573_ _1581_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2733__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4488_ _1508_ _1510_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3508_ _0529_ _0597_ _0524_ _0609_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3439_ _2013_ _0536_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4238__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4705__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4410__A1 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2575__I1 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 net30 X[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 X[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4477__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4229__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3204__I _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2810_ _2075_ _2138_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3790_ _0860_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2741_ _1832_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2963__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _1444_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2672_ Control_Unit.C\[8\] _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4342_ _1373_ _1376_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4273_ _1322_ _1320_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3224_ Control_Unit.T\[14\] _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
.ends

